* Spice description of inverting_mux
* Spice driver version -1217867207
* Date ( dd/mm/yyyy hh:mm:ss ): 10/11/2020 at 14:59:12

* INTERF a0 a1 s sb vdd vss y 


.subckt inverting_mux 1 10 38 20 63 96 87 
* NET 1 = a0
* NET 10 = a1
* NET 20 = sb
* NET 38 = s
* NET 63 = vdd
* NET 87 = y
* NET 96 = vss
Mtr_00008 58 31 90 63 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00007 58 16 62 63 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00006 55 44 88 63 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00005 55 7 61 63 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00004 106 39 82 96 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 106 14 99 96 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 109 19 77 96 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 109 5 97 96 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R11_1 3 2 0.001
R11_2 1 6 0.7
C11_21 1 96 2.17e-15
C11_22 6 96 2.17e-15
R11_3 2 1 0.1
C11_31 2 96 4.2e-16
C11_32 1 96 4.2e-16
R11_4 4 2 0.6
C11_41 4 96 1.75e-15
C11_42 2 96 1.75e-15
R11_5 3 7 450
C11_51 3 96 1.425e-15
C11_52 7 96 1.425e-15
R11_6 5 3 500
C11_61 5 96 1.575e-15
C11_62 3 96 1.575e-15
R10_1 12 11 0.001
R10_2 10 15 0.7
C10_21 10 96 2.17e-15
C10_22 15 96 2.17e-15
R10_3 11 10 0.1
C10_31 11 96 4.2e-16
C10_32 10 96 4.2e-16
R10_4 13 11 0.6
C10_41 13 96 1.75e-15
C10_42 11 96 1.75e-15
R10_5 12 16 450
C10_51 12 96 1.425e-15
C10_52 16 96 1.425e-15
R10_6 14 12 500
C10_61 14 96 1.575e-15
C10_62 12 96 1.575e-15
R9_1 23 22 0.001
R9_2 22 24 0.001
R9_3 24 25 0.001
R9_4 27 26 0.001
R9_5 29 28 0.001
R9_6 35 34 0.001
R9_7 31 35 350
C9_71 31 96 1.125e-15
C9_72 35 96 1.125e-15
R9_8 32 34 0.5
C9_81 32 96 5.75e-16
C9_82 34 96 5.75e-16
R9_9 32 33 0.2
C9_91 32 96 2.875e-16
C9_92 33 96 2.875e-16
R9_10 28 32 0.4
C9_101 28 96 4.6e-16
C9_102 32 96 4.6e-16
R9_11 30 28 0.5
C9_111 30 96 6.325e-16
C9_112 28 96 6.325e-16
R9_12 26 29 0.5
C9_121 26 96 2.4e-15
C9_122 29 96 2.4e-15
R9_13 25 27 0.35
C9_131 25 96 1.8e-15
C9_132 27 96 1.8e-15
R9_14 20 22 0.5
C9_141 20 96 5.75e-16
C9_142 22 96 5.75e-16
R9_15 21 20 0.5
C9_151 21 96 6.325e-16
C9_152 20 96 6.325e-16
R9_16 19 23 400
C9_161 19 96 1.275e-15
C9_162 23 96 1.275e-15
R8_1 49 52 0.001
R8_2 46 45 0.001
R8_3 48 47 0.001
R8_4 41 40 0.001
R8_5 40 42 0.001
R8_6 42 43 0.001
R8_7 39 43 400
C8_71 39 96 1.275e-15
C8_72 43 96 1.275e-15
R8_8 38 42 1
C8_81 38 96 1.15e-15
C8_82 42 96 1.15e-15
R8_9 41 47 0.25
C8_91 41 96 1.2e-15
C8_92 47 96 1.2e-15
R8_10 46 48 0.5
C8_101 46 96 2.4e-15
C8_102 48 96 2.4e-15
R8_11 50 51 0.2
C8_111 50 96 2.875e-16
C8_112 51 96 2.875e-16
R8_12 45 50 0.9
C8_121 45 96 1.035e-15
C8_122 50 96 1.035e-15
R8_13 50 52 0.5
C8_131 50 96 5.75e-16
C8_132 52 96 5.75e-16
R8_14 44 49 350
C8_141 44 96 1.125e-15
C8_142 49 96 1.125e-15
R5_1 62 68 0.001
R5_2 73 72 0.001
R5_3 61 63 0.001
R5_4 67 66 0.001
R5_5 66 69 0.001
C5_51 66 96 8.4e-16
C5_52 69 96 8.4e-16
R5_6 65 66 0.1
C5_61 65 96 1.44e-15
C5_62 66 96 1.44e-15
R5_7 63 65 0.1
C5_71 63 96 1.44e-15
C5_72 65 96 1.44e-15
R5_8 64 63 0.001
C5_81 64 96 1.08e-15
C5_82 63 96 1.08e-15
R5_9 72 74 0.001
C5_91 72 96 1.08e-15
C5_92 74 96 1.08e-15
R5_10 71 72 0.1
C5_101 71 96 1.44e-15
C5_102 72 96 1.44e-15
R5_11 68 71 0.1
C5_111 68 96 1.44e-15
C5_112 71 96 1.44e-15
R5_12 70 68 0.001
C5_121 70 96 8.4e-16
C5_122 68 96 8.4e-16
R5_13 69 70 0.001
C5_131 69 96 2.4e-16
C5_132 70 96 2.4e-16
R4_1 77 78 0.001
R4_2 80 79 0.001
R4_3 88 89 0.001
R4_4 84 83 0.001
R4_5 90 91 0.001
R4_6 82 85 0.001
R4_7 85 86 0.1
C4_71 85 96 1.725e-16
C4_72 86 96 1.725e-16
R4_8 91 93 0.1
C4_81 91 96 1.725e-16
C4_82 93 96 1.725e-16
R4_9 87 91 1.1
C4_91 87 96 1.265e-15
C4_92 91 96 1.265e-15
R4_10 83 87 0.5
C4_101 83 96 5.75e-16
C4_102 87 96 5.75e-16
R4_11 86 83 0.2
C4_111 86 96 2.875e-16
C4_112 83 96 2.875e-16
R4_12 80 84 0.5
C4_121 80 96 2.4e-15
C4_122 84 96 2.4e-15
R4_13 89 92 0.1
C4_131 89 96 1.725e-16
C4_132 92 96 1.725e-16
R4_14 79 89 1.6
C4_141 79 96 1.84e-15
C4_142 89 96 1.84e-15
R4_15 81 79 0.2
C4_151 81 96 2.875e-16
C4_152 79 96 2.875e-16
R4_16 78 81 0.1
C4_161 78 96 1.725e-16
C4_162 81 96 1.725e-16
R3_1 99 100 0.001
R3_2 97 96 0.001
R3_3 96 101 0.2
C3_31 96 96 3.72e-15
C3_32 101 96 3.72e-15
R3_4 98 96 0.001
C3_41 98 96 1.08e-15
C3_42 96 96 1.08e-15
R3_5 100 103 0.2
C3_51 100 96 3.96e-15
C3_52 103 96 3.96e-15
R3_6 102 100 0.001
C3_61 102 96 8.4e-16
C3_62 100 96 8.4e-16
R3_7 101 102 0.001
C3_71 101 96 2.4e-16
C3_72 102 96 2.4e-16
.ends inverting_mux

