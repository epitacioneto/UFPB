* Spice description of noc
* Spice driver version -1218047431
* Date ( dd/mm/yyyy hh:mm:ss ): 12/11/2020 at 15:35:50

* INTERF phi phi1 phi2 vdd vss vss1 


.subckt noc 176 98 198 233 299 25 
* NET 25 = vss1
* NET 31 = inv6.i
* NET 49 = inv6.nq
* NET 65 = inv8.i
* NET 81 = inv8.nq
* NET 98 = phi1
* NET 117 = inv0.nq
* NET 137 = inv3.nq
* NET 153 = inv2.nq
* NET 176 = phi
* NET 198 = phi2
* NET 233 = vdd
* NET 245 = nor1.nq
* NET 262 = inv1.nq
* NET 299 = vss
Mtr_00026 242 178 253 233 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00025 204 190 242 233 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00024 119 181 209 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 52 33 238 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 68 49 237 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 84 65 236 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 194 81 235 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 28 106 31 233 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00018 239 125 28 233 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00017 100 143 208 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00016 144 159 207 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 160 268 206 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 269 252 205 233 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 245 189 298 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 297 169 245 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 304 172 117 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 4 42 61 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 3 59 77 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 2 75 93 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 1 91 200 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 44 132 5 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 6 114 44 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 303 140 97 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 302 156 137 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 301 265 153 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 300 248 262 299 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
R17_1 2 11 0.001
R17_2 1 7 0.001
R17_3 3 14 0.001
R17_4 4 17 0.001
R17_5 6 21 0.001
R17_6 5 18 0.001
R17_7 23 24 0.2
C17_71 23 299 3.6e-15
C17_72 24 299 3.6e-15
R17_8 22 23 0.001
C17_81 22 299 2.4e-16
C17_82 23 299 2.4e-16
R17_9 21 22 0.001
C17_91 21 299 8.4e-16
C17_92 22 299 8.4e-16
R17_10 18 21 0.2
C17_101 18 299 2.88e-15
C17_102 21 299 2.88e-15
R17_11 19 18 0.001
C17_111 19 299 8.4e-16
C17_112 18 299 8.4e-16
R17_12 20 19 0.001
C17_121 20 299 2.4e-16
C17_122 19 299 2.4e-16
R17_13 17 20 0.001
C17_131 17 299 8.4e-16
C17_132 20 299 8.4e-16
R17_14 15 17 0.1
C17_141 15 299 2.52e-15
C17_142 17 299 2.52e-15
R17_15 16 15 0.001
C17_151 16 299 2.4e-16
C17_152 15 299 2.4e-16
R17_16 14 16 0.001
C17_161 14 299 8.4e-16
C17_162 16 299 8.4e-16
R17_17 12 14 0.1
C17_171 12 299 2.52e-15
C17_172 14 299 2.52e-15
R17_18 7 8 0.001
C17_181 7 299 8.4e-16
C17_182 8 299 8.4e-16
R17_19 10 7 0.1
C17_191 10 299 2.76e-15
C17_192 7 299 2.76e-15
R17_20 13 12 0.001
C17_201 13 299 2.4e-16
C17_202 12 299 2.4e-16
R17_21 11 13 0.001
C17_211 11 299 8.4e-16
C17_212 13 299 8.4e-16
R17_22 11 25 0.001
C17_221 11 299 7.2e-16
C17_222 25 299 7.2e-16
R17_23 9 25 0.1
C17_231 9 299 1.8e-15
C17_232 25 299 1.8e-15
R17_24 8 9 0.001
C17_241 8 299 2.4e-16
C17_242 9 299 2.4e-16
R15_1 41 40 0.001
R15_2 37 36 0.001
R15_3 39 38 0.001
R15_4 38 31 0.001
R15_5 31 35 0.001
R15_6 31 32 0.001
R15_7 44 45 0.001
R15_8 45 46 0.2
C15_81 45 299 7e-16
C15_82 46 299 7e-16
R15_9 38 46 1
C15_91 38 299 2.8e-15
C15_92 46 299 2.8e-15
R15_10 35 38 0.2
C15_101 35 299 7e-16
C15_102 38 299 7e-16
R15_11 32 35 0.2
C15_111 32 299 7e-16
C15_112 35 299 7e-16
R15_12 37 39 0.5
C15_121 37 299 2.4e-15
C15_122 39 299 2.4e-15
R15_13 40 43 0.5
C15_131 40 299 1.47e-15
C15_132 43 299 1.47e-15
R15_14 36 40 0.5
C15_141 36 299 1.4e-15
C15_142 40 299 1.4e-15
R15_15 34 36 0.5
C15_151 34 299 1.47e-15
C15_152 36 299 1.47e-15
R15_16 41 42 500
C15_161 41 299 1.5e-15
C15_162 42 299 1.5e-15
R15_17 33 41 600
C15_171 33 299 1.875e-15
C15_172 41 299 1.875e-15
R14_1 52 53 0.001
R14_2 52 56 0.001
R14_3 61 62 0.001
R14_4 55 54 0.001
R14_5 51 50 0.001
R14_6 58 57 0.001
R14_7 58 59 500
C14_71 58 299 1.5e-15
C14_72 59 299 1.5e-15
R14_8 49 58 600
C14_81 49 299 1.875e-15
C14_82 58 299 1.875e-15
R14_9 57 60 0.5
C14_91 57 299 1.47e-15
C14_92 60 299 1.47e-15
R14_10 50 57 1
C14_101 50 299 2.8e-15
C14_102 57 299 2.8e-15
R14_11 51 55 0.25
C14_111 51 299 1.2e-15
C14_112 55 299 1.2e-15
R14_12 56 62 1
C14_121 56 299 2.8e-15
C14_122 62 299 2.8e-15
R14_13 53 56 0.2
C14_131 53 299 7e-16
C14_132 56 299 7e-16
R14_14 54 53 0.2
C14_141 54 299 7e-16
C14_142 53 299 7e-16
R13_1 74 73 0.001
R13_2 67 66 0.001
R13_3 70 69 0.001
R13_4 77 78 0.001
R13_5 68 71 0.001
R13_6 68 72 0.001
R13_7 72 78 1
C13_71 72 299 2.8e-15
C13_72 78 299 2.8e-15
R13_8 71 72 0.2
C13_81 71 299 7e-16
C13_82 72 299 7e-16
R13_9 69 71 0.2
C13_91 69 299 7e-16
C13_92 71 299 7e-16
R13_10 67 70 0.25
C13_101 67 299 1.2e-15
C13_102 70 299 1.2e-15
R13_11 73 76 0.5
C13_111 73 299 1.47e-15
C13_112 76 299 1.47e-15
R13_12 66 73 1
C13_121 66 299 2.8e-15
C13_122 73 299 2.8e-15
R13_13 74 75 500
C13_131 74 299 1.5e-15
C13_132 75 299 1.5e-15
R13_14 65 74 600
C13_141 65 299 1.875e-15
C13_142 74 299 1.875e-15
R12_1 84 85 0.001
R12_2 84 88 0.001
R12_3 93 94 0.001
R12_4 87 86 0.001
R12_5 83 82 0.001
R12_6 90 89 0.001
R12_7 90 91 500
C12_71 90 299 1.5e-15
C12_72 91 299 1.5e-15
R12_8 81 90 600
C12_81 81 299 1.875e-15
C12_82 90 299 1.875e-15
R12_9 89 92 0.5
C12_91 89 299 1.47e-15
C12_92 92 299 1.47e-15
R12_10 82 89 1
C12_101 82 299 2.8e-15
C12_102 89 299 2.8e-15
R12_11 83 87 0.25
C12_111 83 299 1.2e-15
C12_112 87 299 1.2e-15
R12_12 88 94 1
C12_121 88 299 2.8e-15
C12_122 94 299 2.8e-15
R12_13 85 88 0.2
C12_131 85 299 7e-16
C12_132 88 299 7e-16
R12_14 86 85 0.2
C12_141 86 299 7e-16
C12_142 85 299 7e-16
R11_1 97 99 0.001
R11_2 100 101 0.001
R11_3 104 103 0.001
R11_4 100 102 0.001
R11_5 104 105 0.001
R11_6 110 109 0.001
R11_7 108 107 0.001
R11_8 106 111 0.001
R11_9 112 114 700
C11_91 112 299 2.1e-15
C11_92 114 299 2.1e-15
R11_10 106 112 150
C11_101 106 299 4.5e-16
C11_102 112 299 4.5e-16
R11_11 111 113 0.5
C11_111 111 299 1.47e-15
C11_112 113 299 1.47e-15
R11_12 107 111 0.7
C11_121 107 299 2.1e-15
C11_122 111 299 2.1e-15
R11_13 108 109 0.1
C11_131 108 299 6e-16
C11_132 109 299 6e-16
R11_14 105 110 0.5
C11_141 105 299 2.4e-15
C11_142 110 299 2.4e-15
R11_15 101 103 0.2
C11_151 101 299 7e-16
C11_152 103 299 7e-16
R11_16 102 101 0.2
C11_161 102 299 7e-16
C11_162 101 299 7e-16
R11_17 98 102 0.5
C11_171 98 299 1.4e-15
C11_172 102 299 1.4e-15
R11_18 99 98 0.5
C11_181 99 299 1.4e-15
C11_182 98 299 1.4e-15
R10_1 117 118 0.001
R10_2 119 120 0.001
R10_3 123 122 0.001
R10_4 119 121 0.001
R10_5 123 124 0.001
R10_6 130 129 0.001
R10_7 127 126 0.001
R10_8 131 133 0.001
R10_9 131 132 500
C10_91 131 299 1.5e-15
C10_92 132 299 1.5e-15
R10_10 125 131 850
C10_101 125 299 2.625e-15
C10_102 131 299 2.625e-15
R10_11 133 134 0.5
C10_111 133 299 1.47e-15
C10_112 134 299 1.47e-15
R10_12 126 133 0.7
C10_121 126 299 2.1e-15
C10_122 133 299 2.1e-15
R10_13 128 126 0.2
C10_131 128 299 7.7e-16
C10_132 126 299 7.7e-16
R10_14 127 129 0.6
C10_141 127 299 3e-15
C10_142 129 299 3e-15
R10_15 124 130 0.6
C10_151 124 299 3e-15
C10_152 130 299 3e-15
R10_16 120 122 0.2
C10_161 120 299 7e-16
C10_162 122 299 7e-16
R10_17 121 120 0.2
C10_171 121 299 7e-16
C10_172 120 299 7e-16
R10_18 118 121 1
C10_181 118 299 2.8e-15
C10_182 121 299 2.8e-15
R9_1 137 138 0.001
R9_2 144 145 0.001
R9_3 148 147 0.001
R9_4 144 146 0.001
R9_5 150 149 0.001
R9_6 142 141 0.001
R9_7 142 143 600
C9_71 142 299 1.875e-15
C9_72 143 299 1.875e-15
R9_8 140 142 500
C9_81 140 299 1.5e-15
C9_82 142 299 1.5e-15
R9_9 141 149 1
C9_91 141 299 2.8e-15
C9_92 149 299 2.8e-15
R9_10 139 141 0.5
C9_101 139 299 1.47e-15
C9_102 141 299 1.47e-15
R9_11 148 150 0.25
C9_111 148 299 1.2e-15
C9_112 150 299 1.2e-15
R9_12 145 147 0.2
C9_121 145 299 7e-16
C9_122 147 299 7e-16
R9_13 146 145 0.2
C9_131 146 299 7e-16
C9_132 145 299 7e-16
R9_14 138 146 1
C9_141 138 299 2.8e-15
C9_142 146 299 2.8e-15
R8_1 153 154 0.001
R8_2 160 161 0.001
R8_3 164 163 0.001
R8_4 160 162 0.001
R8_5 166 165 0.001
R8_6 158 157 0.001
R8_7 158 159 600
C8_71 158 299 1.875e-15
C8_72 159 299 1.875e-15
R8_8 156 158 500
C8_81 156 299 1.5e-15
C8_82 158 299 1.5e-15
R8_9 157 165 1
C8_91 157 299 2.8e-15
C8_92 165 299 2.8e-15
R8_10 155 157 0.5
C8_101 155 299 1.47e-15
C8_102 157 299 1.47e-15
R8_11 164 166 0.25
C8_111 164 299 1.2e-15
C8_112 166 299 1.2e-15
R8_12 161 163 0.2
C8_121 161 299 7e-16
C8_122 163 299 7e-16
R8_13 162 161 0.2
C8_131 162 299 7e-16
C8_132 161 299 7e-16
R8_14 154 162 1
C8_141 154 299 2.8e-15
C8_142 162 299 2.8e-15
R7_1 178 179 0.001
R7_2 171 170 0.001
R7_3 174 173 0.001
R7_4 177 176 0.001
R7_5 177 181 600
C7_51 177 299 1.875e-15
C7_52 181 299 1.875e-15
R7_6 172 177 500
C7_61 172 299 1.5e-15
C7_62 177 299 1.5e-15
R7_7 176 183 1
C7_71 176 299 2.87e-15
C7_72 183 299 2.87e-15
R7_8 173 176 0.2
C7_81 173 299 7e-16
C7_82 176 299 7e-16
R7_9 175 173 0.2
C7_91 175 299 7.7e-16
C7_92 173 299 7.7e-16
R7_10 171 174 1.85
C7_101 171 299 9e-15
C7_102 174 299 9e-15
R7_11 179 182 0.7
C7_111 179 299 2.17e-15
C7_112 182 299 2.17e-15
R7_12 170 179 0.5
C7_121 170 299 1.4e-15
C7_122 179 299 1.4e-15
R7_13 178 180 150
C7_131 178 299 4.5e-16
C7_132 180 299 4.5e-16
R7_14 169 180 700
C7_141 169 299 2.1e-15
C7_142 180 299 2.1e-15
R6_1 187 186 0.001
R6_2 192 191 0.001
R6_3 192 193 0.001
R6_4 196 195 0.001
R6_5 195 197 0.001
R6_6 200 201 0.001
R6_7 194 198 0.001
R6_8 194 199 0.001
R6_9 199 201 1
C6_91 199 299 2.8e-15
C6_92 201 299 2.8e-15
R6_10 198 199 0.2
C6_101 198 299 7e-16
C6_102 199 299 7e-16
R6_11 197 198 0.2
C6_111 197 299 7e-16
C6_112 198 299 7e-16
R6_12 193 196 0.5
C6_121 193 299 2.4e-15
C6_122 196 299 2.4e-15
R6_13 186 191 1
C6_131 186 299 2.8e-15
C6_132 191 299 2.8e-15
R6_14 188 186 0.5
C6_141 188 299 1.47e-15
C6_142 186 299 1.47e-15
R6_15 189 187 500
C6_151 189 299 1.5e-15
C6_152 187 299 1.5e-15
R6_16 187 190 850
C6_161 187 299 2.625e-15
C6_162 190 299 2.625e-15
R5_1 205 214 0.001
R5_2 237 218 0.001
R5_3 206 218 0.001
R5_4 236 214 0.001
R5_5 204 210 0.001
R5_6 238 221 0.001
R5_7 207 221 0.001
R5_8 235 232 0.001
R5_9 239 234 0.001
R5_10 208 226 0.001
R5_11 209 227 0.001
R5_12 230 231 0.001
C5_121 230 299 2.145e-15
C5_122 231 299 2.145e-15
R5_13 227 230 0.001
C5_131 227 299 2.34e-15
C5_132 230 299 2.34e-15
R5_14 228 227 0.001
C5_141 228 299 1.365e-15
C5_142 227 299 1.365e-15
R5_15 229 228 0.001
C5_151 229 299 3.9e-16
C5_152 228 299 3.9e-16
R5_16 225 229 0.001
C5_161 225 299 1.755e-15
C5_162 229 299 1.755e-15
R5_17 226 225 0.001
C5_171 226 299 2.34e-15
C5_172 225 299 2.34e-15
R5_18 223 226 0.001
C5_181 223 299 1.365e-15
C5_182 226 299 1.365e-15
R5_19 224 223 0.001
C5_191 224 299 3.9e-16
C5_192 223 299 3.9e-16
R5_20 224 234 0.001
C5_201 224 299 5.85e-16
C5_202 234 299 5.85e-16
R5_21 222 234 0.001
C5_211 222 299 1.17e-15
C5_212 234 299 1.17e-15
R5_22 221 222 0.001
C5_221 221 299 1.95e-15
C5_222 222 299 1.95e-15
R5_23 220 221 0.001
C5_231 220 299 1.95e-15
C5_232 221 299 1.95e-15
R5_24 212 232 0.001
C5_241 212 299 1.365e-15
C5_242 232 299 1.365e-15
R5_25 210 232 0.001
C5_251 210 299 2.73e-15
C5_252 232 299 2.73e-15
R5_26 211 210 0.001
C5_261 211 299 1.755e-15
C5_262 210 299 1.755e-15
R5_27 214 216 0.001
C5_271 214 299 1.95e-15
C5_272 216 299 1.95e-15
R5_28 213 215 0.001
C5_281 213 299 1.755e-15
C5_282 215 299 1.755e-15
R5_29 212 213 0.001
C5_291 212 299 3.9e-16
C5_292 213 299 3.9e-16
R5_30 219 220 0.001
C5_301 219 299 1.95e-15
C5_302 220 299 1.95e-15
R5_31 218 219 0.001
C5_311 218 299 1.95e-15
C5_312 219 299 1.95e-15
R5_32 217 218 0.001
C5_321 217 299 1.95e-15
C5_322 218 299 1.95e-15
R5_33 216 217 0.001
C5_331 216 299 1.95e-15
C5_332 217 299 1.95e-15
R5_34 216 233 0.001
C5_341 216 299 4.8e-16
C5_342 233 299 4.8e-16
R5_35 214 233 0.001
C5_351 214 299 7.2e-16
C5_352 233 299 7.2e-16
R5_36 215 214 0.001
C5_361 215 299 1.95e-15
C5_362 214 299 1.95e-15
R3_1 245 246 0.001
R3_2 253 255 0.001
R3_3 253 256 0.001
R3_4 257 256 0.001
R3_5 253 254 0.001
R3_6 259 258 0.001
R3_7 250 251 0.001
R3_8 250 252 600
C3_81 250 299 1.875e-15
C3_82 252 299 1.875e-15
R3_9 248 250 500
C3_91 248 299 1.5e-15
C3_92 250 299 1.5e-15
R3_10 251 258 1
C3_101 251 299 2.8e-15
C3_102 258 299 2.8e-15
R3_11 249 251 0.5
C3_111 249 299 1.47e-15
C3_112 251 299 1.47e-15
R3_12 257 259 0.25
C3_121 257 299 1.2e-15
C3_122 259 299 1.2e-15
R3_13 255 256 0.2
C3_131 255 299 7e-16
C3_132 256 299 7e-16
R3_14 254 255 0.2
C3_141 254 299 7e-16
C3_142 255 299 7e-16
R3_15 247 254 1
C3_151 247 299 2.8e-15
C3_152 254 299 2.8e-15
R3_16 246 247 0.2
C3_161 246 299 7e-16
C3_162 247 299 7e-16
R2_1 262 263 0.001
R2_2 270 269 0.001
R2_3 273 272 0.001
R2_4 271 269 0.001
R2_5 275 274 0.001
R2_6 267 266 0.001
R2_7 267 268 600
C2_71 267 299 1.875e-15
C2_72 268 299 1.875e-15
R2_8 265 267 500
C2_81 265 299 1.5e-15
C2_82 267 299 1.5e-15
R2_9 266 274 1
C2_91 266 299 2.8e-15
C2_92 274 299 2.8e-15
R2_10 264 266 0.5
C2_101 264 299 1.47e-15
C2_102 266 299 1.47e-15
R2_11 272 275 0.25
C2_111 272 299 1.2e-15
C2_112 275 299 1.2e-15
R2_12 270 273 0.2
C2_121 270 299 7e-16
C2_122 273 299 7e-16
R2_13 271 270 0.2
C2_131 271 299 7e-16
C2_132 270 299 7e-16
R2_14 263 271 1
C2_141 263 299 2.8e-15
C2_142 271 299 2.8e-15
R1_1 297 278 0.001
R1_2 298 279 0.001
R1_3 300 281 0.001
R1_4 301 284 0.001
R1_5 302 287 0.001
R1_6 303 290 0.001
R1_7 304 294 0.001
R1_8 294 296 0.1
C1_81 294 299 2.76e-15
C1_82 296 299 2.76e-15
R1_9 295 294 0.001
C1_91 295 299 8.4e-16
C1_92 294 299 8.4e-16
R1_10 291 295 0.001
C1_101 291 299 2.4e-16
C1_102 295 299 2.4e-16
R1_11 290 291 0.1
C1_111 290 299 2.52e-15
C1_112 291 299 2.52e-15
R1_12 292 290 0.001
C1_121 292 299 8.4e-16
C1_122 290 299 8.4e-16
R1_13 293 292 0.001
C1_131 293 299 2.4e-16
C1_132 292 299 2.4e-16
R1_14 287 293 0.1
C1_141 287 299 2.52e-15
C1_142 293 299 2.52e-15
R1_15 288 287 0.001
C1_151 288 299 8.4e-16
C1_152 287 299 8.4e-16
R1_16 289 288 0.001
C1_161 289 299 2.4e-16
C1_162 288 299 2.4e-16
R1_17 284 289 0.1
C1_171 284 299 2.52e-15
C1_172 289 299 2.52e-15
R1_18 285 284 0.001
C1_181 285 299 8.4e-16
C1_182 284 299 8.4e-16
R1_19 286 285 0.001
C1_191 286 299 2.4e-16
C1_192 285 299 2.4e-16
R1_20 299 286 0.1
C1_201 299 299 1.56e-15
C1_202 286 299 1.56e-15
R1_21 281 299 0.001
C1_211 281 299 9.6e-16
C1_212 299 299 9.6e-16
R1_22 282 281 0.001
C1_221 282 299 8.4e-16
C1_222 281 299 8.4e-16
R1_23 283 282 0.001
C1_231 283 299 2.4e-16
C1_232 282 299 2.4e-16
R1_24 278 283 0.001
C1_241 278 299 8.4e-16
C1_242 283 299 8.4e-16
R1_25 279 278 0.2
C1_251 279 299 2.88e-15
C1_252 278 299 2.88e-15
R1_26 280 279 0.001
C1_261 280 299 1.08e-15
C1_262 279 299 1.08e-15
.ends noc

