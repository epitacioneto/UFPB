* Spice description of ff_m_e_noc_roteado
* Spice driver version -1217539527
* Date ( dd/mm/yyyy hh:mm:ss ): 19/11/2020 at 16:17:05

* INTERF a ck phi_1 phi_2 q vdd vss 


.subckt ff_m_e_noc_roteado 29 22 14 30 12 34 21 
* NET 1 = nock.i9
* NET 2 = nock.i7
* NET 3 = nock.i8
* NET 4 = nock.ck_b
* NET 6 = nock.i6
* NET 9 = nock.i3
* NET 10 = ff.la_e.q_b
* NET 11 = nock.i4
* NET 12 = q
* NET 13 = ff.la_e.b
* NET 14 = phi_1
* NET 21 = vss
* NET 22 = ck
* NET 23 = nock.i2
* NET 25 = nock.i1
* NET 26 = ff.la_m.q_b
* NET 27 = ff.q_m
* NET 28 = ff.la_m.b
* NET 29 = a
* NET 30 = phi_2
* NET 34 = vdd
Mtr_00058 34 33 27 34 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00057 35 29 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 31 30 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 32 30 33 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 33 31 35 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 34 28 32 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 26 27 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 28 26 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 23 25 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 24 30 25 34 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00048 34 22 24 34 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00047 34 17 12 34 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00046 8 27 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00045 15 14 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 7 14 17 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 17 15 8 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 34 13 7 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 14 11 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 11 9 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 13 10 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 9 23 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 10 12 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 5 14 6 34 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00035 34 4 5 34 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00034 3 2 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 2 6 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00032 30 1 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 4 22 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 1 3 34 34 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00029 21 29 20 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 20 30 33 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 21 30 31 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00026 33 31 19 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00025 19 28 21 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00024 27 33 21 21 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 21 27 26 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 21 26 28 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00021 21 25 23 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00020 25 22 21 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 21 30 25 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 21 27 18 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00017 18 14 17 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00016 21 14 15 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00015 17 15 16 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00014 16 13 21 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00013 12 17 21 21 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 21 11 14 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 21 9 11 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 21 10 13 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 21 23 9 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 21 12 10 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 6 4 21 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 21 14 6 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 21 2 3 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 21 6 2 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 21 1 30 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 21 22 4 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 21 3 1 21 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C36 1 21 5.497e-14
C35 2 21 5.257e-14
C34 3 21 6.457e-14
C33 4 21 6.722e-14
C31 6 21 6.081e-14
C27 9 21 5.377e-14
C26 10 21 5.377e-14
C25 11 21 5.017e-14
C24 12 21 6.541e-14
C23 13 21 6.328e-14
C22 14 21 9.798e-14
C21 15 21 2.356e-14
C19 17 21 1.932e-14
C15 21 21 4.43001e-13
C14 22 21 7.483e-14
C13 23 21 5.449e-14
C11 25 21 5.121e-14
C10 26 21 5.017e-14
C9 27 21 9.346e-14
C8 28 21 6.208e-14
C7 29 21 3.309e-14
C6 30 21 1.2798e-13
C5 31 21 2.356e-14
C3 33 21 1.932e-14
C2 34 21 4.71001e-13
.ends ff_m_e_noc_roteado

