* Spice description of inv3_s
* Spice driver version -1217543623
* Date ( dd/mm/yyyy hh:mm:ss ): 17/10/2020 at 21:44:16

* INTERF a vdd vss y1 y2 y3 


.subckt inv3_s 9 33 69 47 83 5 
* NET 5 = y3
* NET 9 = a
* NET 33 = vdd
* NET 47 = y1
* NET 69 = vss
* NET 83 = y2
Mtr_00006 4 85 20 33 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 84 49 19 33 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 48 15 18 33 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 1 75 62 69 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 72 39 57 69 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 36 13 54 69 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R6_1 1 2 0.001
R6_2 4 5 0.001
R6_3 5 6 0.4
C6_31 5 69 1.365e-15
C6_32 6 69 1.365e-15
R6_4 2 5 0.9
C6_41 2 69 2.765e-15
C6_42 5 69 2.765e-15
R6_5 3 2 0.001
C6_51 3 69 2.1e-16
C6_52 2 69 2.1e-16
R5_1 11 10 0.001
R5_2 9 14 0.7
C5_21 9 69 2.17e-15
C5_22 14 69 2.17e-15
R5_3 10 9 0.1
C5_31 10 69 4.2e-16
C5_32 9 69 4.2e-16
R5_4 12 10 0.6
C5_41 12 69 1.75e-15
C5_42 10 69 1.75e-15
R5_5 11 15 550
C5_51 11 69 1.65e-15
C5_52 15 69 1.65e-15
R5_6 13 11 500
C5_61 13 69 1.575e-15
C5_62 11 69 1.575e-15
R4_1 18 21 0.001
R4_2 19 26 0.001
R4_3 20 28 0.001
R4_4 31 32 0.001
C4_41 31 69 1.32e-15
C4_42 32 69 1.32e-15
R4_5 28 31 0.1
C4_51 28 69 1.44e-15
C4_52 31 69 1.44e-15
R4_6 29 28 0.001
C4_61 29 69 8.4e-16
C4_62 28 69 8.4e-16
R4_7 30 29 0.001
C4_71 30 69 2.4e-16
C4_72 29 69 2.4e-16
R4_8 27 30 0.001
C4_81 27 69 1.08e-15
C4_82 30 69 1.08e-15
R4_9 26 27 0.1
C4_91 26 69 1.44e-15
C4_92 27 69 1.44e-15
R4_10 24 26 0.001
C4_101 24 69 8.4e-16
C4_102 26 69 8.4e-16
R4_11 25 24 0.001
C4_111 25 69 2.4e-16
C4_112 24 69 2.4e-16
R4_12 23 25 0.001
C4_121 23 69 1.08e-15
C4_122 25 69 1.08e-15
R4_13 23 33 0.001
C4_131 23 69 7.2e-16
C4_132 33 69 7.2e-16
R4_14 21 33 0.001
C4_141 21 69 7.2e-16
C4_142 33 69 7.2e-16
R4_15 22 21 0.001
C4_151 22 69 1.08e-15
C4_152 21 69 1.08e-15
R3_1 36 37 0.001
R3_2 48 47 0.001
R3_3 42 41 0.001
R3_4 45 44 0.001
R3_5 43 46 0.001
R3_6 43 49 550
C3_61 43 69 1.65e-15
C3_62 49 69 1.65e-15
R3_7 39 43 500
C3_71 39 69 1.575e-15
C3_72 43 69 1.575e-15
R3_8 44 51 0.7
C3_81 44 69 2.17e-15
C3_82 51 69 2.17e-15
R3_9 46 44 0.1
C3_91 46 69 4.2e-16
C3_92 44 69 4.2e-16
R3_10 40 46 0.6
C3_101 40 69 1.75e-15
C3_102 46 69 1.75e-15
R3_11 42 45 0.25
C3_111 42 69 1.2e-15
C3_112 45 69 1.2e-15
R3_12 47 50 0.4
C3_121 47 69 1.365e-15
C3_122 50 69 1.365e-15
R3_13 41 47 0.2
C3_131 41 69 8.05e-16
C3_132 47 69 8.05e-16
R3_14 37 41 0.7
C3_141 37 69 1.96e-15
C3_142 41 69 1.96e-15
R3_15 38 37 0.001
C3_151 38 69 2.1e-16
C3_152 37 69 2.1e-16
R2_1 57 61 0.001
R2_2 54 55 0.001
R2_3 62 64 0.001
R2_4 67 68 0.001
C2_41 67 69 6e-16
C2_42 68 69 6e-16
R2_5 64 67 0.1
C2_51 64 69 2.16e-15
C2_52 67 69 2.16e-15
R2_6 65 64 0.001
C2_61 65 69 8.4e-16
C2_62 64 69 8.4e-16
R2_7 58 59 0.001
C2_71 58 69 3.6e-16
C2_72 59 69 3.6e-16
R2_8 58 69 0.001
C2_81 58 69 1.2e-15
C2_82 69 69 1.2e-15
R2_9 55 69 0.001
C2_91 55 69 9.6e-16
C2_92 69 69 9.6e-16
R2_10 56 55 0.001
C2_101 56 69 1.08e-15
C2_102 55 69 1.08e-15
R2_11 66 65 0.001
C2_111 66 69 2.4e-16
C2_112 65 69 2.4e-16
R2_12 63 66 0.001
C2_121 63 69 3.6e-16
C2_122 66 69 3.6e-16
R2_13 61 63 0.1
C2_131 61 69 2.16e-15
C2_132 63 69 2.16e-15
R2_14 60 61 0.001
C2_141 60 69 8.4e-16
C2_142 61 69 8.4e-16
R2_15 59 60 0.001
C2_151 59 69 2.4e-16
C2_152 60 69 2.4e-16
R1_1 72 73 0.001
R1_2 84 83 0.001
R1_3 78 77 0.001
R1_4 81 80 0.001
R1_5 79 82 0.001
R1_6 79 85 550
C1_61 79 69 1.65e-15
C1_62 85 69 1.65e-15
R1_7 75 79 500
C1_71 75 69 1.575e-15
C1_72 79 69 1.575e-15
R1_8 80 87 0.7
C1_81 80 69 2.17e-15
C1_82 87 69 2.17e-15
R1_9 82 80 0.1
C1_91 82 69 4.2e-16
C1_92 80 69 4.2e-16
R1_10 76 82 0.6
C1_101 76 69 1.75e-15
C1_102 82 69 1.75e-15
R1_11 78 81 0.25
C1_111 78 69 1.2e-15
C1_112 81 69 1.2e-15
R1_12 83 86 0.4
C1_121 83 69 1.365e-15
C1_122 86 69 1.365e-15
R1_13 77 83 0.2
C1_131 77 69 8.05e-16
C1_132 83 69 8.05e-16
R1_14 73 77 0.7
C1_141 73 69 1.96e-15
C1_142 77 69 1.96e-15
R1_15 74 73 0.001
C1_151 74 69 2.1e-16
C1_152 73 69 2.1e-16
.ends inv3_s

