* Spice description of tristate_inverter
* Spice driver version -1217633735
* Date ( dd/mm/yyyy hh:mm:ss ):  5/11/2020 at 14:34:43

* INTERF a enable vdd vss y 


.subckt tristate_inverter 13 6 27 60 42 
* NET 6 = enable
* NET 13 = a
* NET 27 = vdd
* NET 42 = y
* NET 60 = vss
Mtr_00006 51 9 25 27 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00005 22 19 26 27 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00004 22 53 43 27 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 48 1 61 60 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 70 17 63 60 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 70 4 38 60 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R8_1 8 7 0.001
R8_2 5 4 250
C8_21 5 60 8.25e-16
C8_22 4 60 8.25e-16
R8_3 6 10 0.7
C8_31 6 60 2.17e-15
C8_32 10 60 2.17e-15
R8_4 7 6 0.1
C8_41 7 60 4.2e-16
C8_42 6 60 4.2e-16
R8_5 2 7 0.6
C8_51 2 60 1.75e-15
C8_52 7 60 1.75e-15
R8_6 3 5 1050
C8_61 3 60 3.15e-15
C8_62 5 60 3.15e-15
R8_7 3 1 250
C8_71 3 60 8.25e-16
C8_72 1 60 8.25e-16
R8_8 8 9 450
C8_81 8 60 1.425e-15
C8_82 9 60 1.425e-15
R8_9 1 8 500
C8_91 1 60 1.575e-15
C8_92 8 60 1.575e-15
R7_1 15 14 0.001
R7_2 13 18 0.7
C7_21 13 60 2.17e-15
C7_22 18 60 2.17e-15
R7_3 14 13 0.1
C7_31 14 60 4.2e-16
C7_32 13 60 4.2e-16
R7_4 16 14 0.6
C7_41 16 60 1.75e-15
C7_42 14 60 1.75e-15
R7_5 15 19 450
C7_51 15 60 1.425e-15
C7_52 19 60 1.425e-15
R7_6 17 15 500
C7_61 17 60 1.575e-15
C7_62 15 60 1.575e-15
R5_1 25 27 0.001
R5_2 34 33 0.001
R5_3 26 31 0.001
R5_4 33 35 0.001
C5_41 33 60 1.08e-15
C5_42 35 60 1.08e-15
R5_5 32 33 0.1
C5_51 32 60 1.44e-15
C5_52 33 60 1.44e-15
R5_6 31 32 0.1
C5_61 31 60 1.44e-15
C5_62 32 60 1.44e-15
R5_7 29 31 0.001
C5_71 29 60 8.4e-16
C5_72 31 60 8.4e-16
R5_8 30 29 0.001
C5_81 30 60 2.4e-16
C5_82 29 60 2.4e-16
R5_9 27 30 0.1
C5_91 27 60 2.52e-15
C5_92 30 60 2.52e-15
R5_10 28 27 0.001
C5_101 28 60 1.08e-15
C5_102 27 60 1.08e-15
R4_1 38 39 0.001
R4_2 43 44 0.001
R4_3 44 45 0.1
C4_31 44 60 1.725e-16
C4_32 45 60 1.725e-16
R4_4 42 44 0.8
C4_41 42 60 9.2e-16
C4_42 44 60 9.2e-16
R4_5 40 42 0.8
C4_51 40 60 9.775e-16
C4_52 42 60 9.775e-16
R4_6 41 40 0.2
C4_61 41 60 2.3e-16
C4_62 40 60 2.3e-16
R4_7 39 41 0.1
C4_71 39 60 1.725e-16
C4_72 41 60 1.725e-16
R3_1 48 49 0.001
R3_2 55 54 0.001
R3_3 51 52 0.001
R3_4 53 56 300
C3_41 53 60 9.75e-16
C3_42 56 60 9.75e-16
R3_5 55 56 900
C3_51 55 60 2.7e-15
C3_52 56 60 2.7e-15
R3_6 54 57 0.1
C3_61 54 60 3.5e-16
C3_62 57 60 3.5e-16
R3_7 52 54 0.3
C3_71 52 60 9.8e-16
C3_72 54 60 9.8e-16
R3_8 49 52 1
C3_81 49 60 2.8e-15
C3_82 52 60 2.8e-15
R3_9 50 49 0.001
C3_91 50 60 2.1e-16
C3_92 49 60 2.1e-16
R2_1 63 64 0.001
R2_2 61 60 0.001
R2_3 60 65 0.1
C2_31 60 60 2.52e-15
C2_32 65 60 2.52e-15
R2_4 62 60 0.001
C2_41 62 60 1.08e-15
C2_42 60 60 1.08e-15
R2_5 64 67 0.2
C2_51 64 60 3.96e-15
C2_52 67 60 3.96e-15
R2_6 66 64 0.001
C2_61 66 60 8.4e-16
C2_62 64 60 8.4e-16
R2_7 65 66 0.001
C2_71 65 60 2.4e-16
C2_72 66 60 2.4e-16
.ends tristate_inverter

