* Spice description of nand2_teste
* Spice driver version -1217895879
* Date ( dd/mm/yyyy hh:mm:ss ):  2/11/2020 at 19:33:27

* INTERF a b vdd vss y 


.subckt nand2_teste 10 4 21 28 41 
* NET 4 = b
* NET 10 = a
* NET 21 = vdd
* NET 28 = vss
* NET 41 = y
Mtr_00004 42 2 20 21 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00003 42 16 19 21 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00002 36 1 39 28 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00001 36 14 29 28 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
R5_1 6 5 0.001
R5_2 3 2 450
C5_21 3 28 1.35e-15
C5_22 2 28 1.35e-15
R5_3 1 3 550
C5_31 1 28 1.65e-15
C5_32 3 28 1.65e-15
R5_4 5 7 0.9
C5_41 5 28 2.59e-15
C5_42 7 28 2.59e-15
R5_5 4 5 0.1
C5_51 4 28 2.8e-16
C5_52 5 28 2.8e-16
R5_6 3 6 200
C5_61 3 28 6e-16
C5_62 6 28 6e-16
R4_1 12 11 0.001
R4_2 11 15 0.9
C4_21 11 28 2.59e-15
C4_22 15 28 2.59e-15
R4_3 10 11 0.1
C4_31 10 28 2.8e-16
C4_32 11 28 2.8e-16
R4_4 13 10 0.5
C4_41 13 28 1.47e-15
C4_42 10 28 1.47e-15
R4_5 12 16 450
C4_51 12 28 1.35e-15
C4_52 16 28 1.35e-15
R4_6 14 12 550
C4_61 14 28 1.65e-15
C4_62 12 28 1.65e-15
R3_1 19 21 0.001
R3_2 20 24 0.001
R3_3 24 25 0.001
C3_31 24 28 1.08e-15
C3_32 25 28 1.08e-15
R3_4 23 24 0.1
C3_41 23 28 1.44e-15
C3_42 24 28 1.44e-15
R3_5 21 23 0.1
C3_51 21 28 1.44e-15
C3_52 23 28 1.44e-15
R3_6 22 21 0.001
C3_61 22 28 1.08e-15
C3_62 21 28 1.08e-15
R2_1 29 28 0.001
R2_2 30 28 0.001
C2_21 30 28 1.08e-15
C2_22 28 28 1.08e-15
R2_3 32 33 0.001
C2_31 32 28 1.2e-15
C2_32 33 28 1.2e-15
R2_4 31 32 0.001
C2_41 31 28 1.32e-15
C2_42 32 28 1.32e-15
R2_5 28 31 0.1
C2_51 28 28 1.44e-15
C2_52 31 28 1.44e-15
R1_1 36 37 0.001
R1_2 39 40 0.001
R1_3 42 43 0.001
R1_4 43 44 0.2
C1_41 43 28 7.7e-16
C1_42 44 28 7.7e-16
R1_5 41 43 0.7
C1_51 41 28 2.1e-15
C1_52 43 28 2.1e-15
R1_6 37 41 0.4
C1_61 37 28 1.26e-15
C1_62 41 28 1.26e-15
R1_7 38 37 0.001
C1_71 38 28 2.1e-16
C1_72 37 28 2.1e-16
R1_8 37 40 0.6
C1_81 37 28 6.9e-16
C1_82 40 28 6.9e-16
.ends nand2_teste

