* Spice description of inversor_gordo
* Spice driver version -1217691079
* Date ( dd/mm/yyyy hh:mm:ss ): 18/10/2020 at 16:19:27

* INTERF a vdd vss y 


.subckt inversor_gordo 1 13 30 19 
* NET 1 = a
* NET 13 = vdd
* NET 19 = y
* NET 30 = vss
Mtr_00002 22 7 10 13 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 18 5 27 30 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
R4_1 3 2 0.001
R4_2 1 6 0.7
C4_21 1 30 2.17e-15
C4_22 6 30 2.17e-15
R4_3 2 1 0.1
C4_31 2 30 4.2e-16
C4_32 1 30 4.2e-16
R4_4 4 2 0.6
C4_41 4 30 1.75e-15
C4_42 2 30 1.75e-15
R4_5 3 7 650
C4_51 3 30 2.025e-15
C4_52 7 30 2.025e-15
R4_6 5 3 550
C4_61 5 30 1.725e-15
C4_62 3 30 1.725e-15
R3_1 10 11 0.001
R3_2 14 15 0.001
C3_21 14 30 1.32e-15
C3_22 15 30 1.32e-15
R3_3 14 13 0.001
C3_31 14 30 7.2e-16
C3_32 13 30 7.2e-16
R3_4 11 13 0.001
C3_41 11 30 7.2e-16
C3_42 13 30 7.2e-16
R3_5 12 11 0.001
C3_51 12 30 1.08e-15
C3_52 11 30 1.08e-15
R2_1 18 20 0.001
R2_2 22 23 0.001
R2_3 23 24 0.4
C2_31 23 30 1.33e-15
C2_32 24 30 1.33e-15
R2_4 19 23 0.8
C2_41 19 30 2.24e-15
C2_42 23 30 2.24e-15
R2_5 20 19 0.2
C2_51 20 30 5.6e-16
C2_52 19 30 5.6e-16
R2_6 21 20 0.001
C2_61 21 30 2.1e-16
C2_62 20 30 2.1e-16
R1_1 27 28 0.001
R1_2 31 32 0.001
C1_21 31 30 6e-16
C1_22 32 30 6e-16
R1_3 31 30 0.001
C1_31 31 30 1.2e-15
C1_32 30 30 1.2e-15
R1_4 28 30 0.001
C1_41 28 30 9.6e-16
C1_42 30 30 9.6e-16
R1_5 29 28 0.001
C1_51 29 30 1.08e-15
C1_52 28 30 1.08e-15
.ends inversor_gordo

