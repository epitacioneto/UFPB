
.include inversor_equilibrado.spi

.model tp pmos level = 54
.model tn nmos level = 54

* a vdd vss y
X1 10 20 30 40 inversor_equilibrado

V1 10 30 pulse(0 1.8 1ns 1ps 1ps 1ns 2ns)
V2 20 30 1.8V
V3 30 0 0V

.tran 0.0001 3ns
.end
