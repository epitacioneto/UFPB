
.include inv3_s.spi

* a vdd vss y1 y2 y3
X1 10 40 30 20 21 22 inv3_s

Vdd 40 30 1.8V
Vss 30 0 0.0V
V1 10 30 pulse(0.716V 1.123V 0 1ps 1ps 4ns 8ns)

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.1n 16n

.end
