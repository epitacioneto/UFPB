* Spice description of fo4_eq2
* Spice driver version -1218260423
* Date ( dd/mm/yyyy hh:mm:ss ): 19/10/2020 at 22:42:07

* INTERF a vdd vss1 vss2 y 


.subckt fo4_eq2 47 77 105 16 127 
* NET 16 = vss2
* NET 47 = a
* NET 77 = vdd
* NET 105 = vss1
* NET 127 = y
Mtr_00012 145 54 76 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 119 50 61 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 19 142 79 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 38 126 63 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 27 141 78 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 85 125 62 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 151 57 1 105 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00005 108 46 90 105 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00004 22 154 3 105 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 35 113 98 105 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 30 153 2 105 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 82 112 93 105 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R9_1 1 4 0.001
R9_2 2 9 0.001
R9_3 3 11 0.001
R9_4 14 15 0.001
C9_41 14 105 6e-16
C9_42 15 105 6e-16
R9_5 11 14 0.1
C9_51 11 105 2.16e-15
C9_52 14 105 2.16e-15
R9_6 12 11 0.001
C9_61 12 105 8.4e-16
C9_62 11 105 8.4e-16
R9_7 13 12 0.001
C9_71 13 105 2.4e-16
C9_72 12 105 2.4e-16
R9_8 10 13 0.001
C9_81 10 105 3.6e-16
C9_82 13 105 3.6e-16
R9_9 10 16 0.1
C9_91 10 105 1.44e-15
C9_92 16 105 1.44e-15
R9_10 9 16 0.001
C9_101 9 105 7.2e-16
C9_102 16 105 7.2e-16
R9_11 7 9 0.001
C9_111 7 105 8.4e-16
C9_112 9 105 8.4e-16
R9_12 8 7 0.001
C9_121 8 105 2.4e-16
C9_122 7 105 2.4e-16
R9_13 6 8 0.001
C9_131 6 105 3.6e-16
C9_132 8 105 3.6e-16
R9_14 4 6 0.1
C9_141 4 105 2.16e-15
C9_142 6 105 2.16e-15
R9_15 5 4 0.001
C9_151 5 105 1.08e-15
C9_152 4 105 1.08e-15
R8_1 22 23 0.001
R8_2 19 20 0.001
R8_3 23 24 0.001
C8_31 23 105 2.1e-16
C8_32 24 105 2.1e-16
R8_4 20 23 1
C8_41 20 105 2.8e-15
C8_42 23 105 2.8e-15
R8_5 21 20 0.4
C8_51 21 105 1.33e-15
C8_52 20 105 1.33e-15
R7_1 30 31 0.001
R7_2 27 28 0.001
R7_3 31 32 0.001
C7_31 31 105 2.1e-16
C7_32 32 105 2.1e-16
R7_4 28 31 1
C7_41 28 105 2.8e-15
C7_42 31 105 2.8e-15
R7_5 29 28 0.4
C7_51 29 105 1.33e-15
C7_52 28 105 1.33e-15
R6_1 35 36 0.001
R6_2 38 39 0.001
R6_3 39 40 0.4
C6_31 39 105 1.33e-15
C6_32 40 105 1.33e-15
R6_4 36 39 1
C6_41 36 105 2.8e-15
C6_42 39 105 2.8e-15
R6_5 37 36 0.001
C6_51 37 105 2.1e-16
C6_52 36 105 2.1e-16
R5_1 44 43 0.001
R5_2 48 47 0.001
R5_3 48 49 0.001
R5_4 52 51 0.001
R5_5 51 53 0.001
R5_6 56 55 0.001
R5_7 56 57 500
C5_71 56 105 1.575e-15
C5_72 57 105 1.575e-15
R5_8 54 56 550
C5_81 54 105 1.65e-15
C5_82 56 105 1.65e-15
R5_9 55 58 0.6
C5_91 55 105 1.75e-15
C5_92 58 105 1.75e-15
R5_10 53 55 0.9
C5_101 53 105 2.52e-15
C5_102 55 105 2.52e-15
R5_11 49 52 0.5
C5_111 49 105 2.4e-15
C5_112 52 105 2.4e-15
R5_12 43 47 0.9
C5_121 43 105 2.52e-15
C5_122 47 105 2.52e-15
R5_13 45 43 0.6
C5_131 45 105 1.75e-15
C5_132 43 105 1.75e-15
R5_14 44 50 550
C5_141 44 105 1.65e-15
C5_142 50 105 1.65e-15
R5_15 46 44 500
C5_151 46 105 1.575e-15
C5_152 44 105 1.575e-15
R4_1 62 67 0.001
R4_2 76 64 0.001
R4_3 78 67 0.001
R4_4 63 73 0.001
R4_5 79 73 0.001
R4_6 61 64 0.001
R4_7 66 77 0.001
C4_71 66 105 7.2e-16
C4_72 77 105 7.2e-16
R4_8 64 77 0.001
C4_81 64 105 7.2e-16
C4_82 77 105 7.2e-16
R4_9 74 75 0.001
C4_91 74 105 2.145e-15
C4_92 75 105 2.145e-15
R4_10 73 74 0.001
C4_101 73 105 2.34e-15
C4_102 74 105 2.34e-15
R4_11 71 73 0.001
C4_111 71 105 1.365e-15
C4_112 73 105 1.365e-15
R4_12 66 68 0.001
C4_121 66 105 1.755e-15
C4_122 68 105 1.755e-15
R4_13 64 66 0.001
C4_131 64 105 2.34e-15
C4_132 66 105 2.34e-15
R4_14 65 64 0.001
C4_141 65 105 1.755e-15
C4_142 64 105 1.755e-15
R4_15 72 71 0.001
C4_151 72 105 3.9e-16
C4_152 71 105 3.9e-16
R4_16 70 72 0.001
C4_161 70 105 1.755e-15
C4_162 72 105 1.755e-15
R4_17 67 70 0.001
C4_171 67 105 2.34e-15
C4_172 70 105 2.34e-15
R4_18 69 67 0.001
C4_181 69 105 1.365e-15
C4_182 67 105 1.365e-15
R4_19 68 69 0.001
C4_191 68 105 3.9e-16
C4_192 69 105 3.9e-16
R3_1 82 83 0.001
R3_2 85 86 0.001
R3_3 86 87 0.4
C3_31 86 105 1.33e-15
C3_32 87 105 1.33e-15
R3_4 83 86 1
C3_41 83 105 2.8e-15
C3_42 86 105 2.8e-15
R3_5 84 83 0.001
C3_51 84 105 2.1e-16
C3_52 83 105 2.1e-16
R2_1 90 91 0.001
R2_2 93 97 0.001
R2_3 98 100 0.001
R2_4 103 104 0.001
C2_41 103 105 6e-16
C2_42 104 105 6e-16
R2_5 100 103 0.1
C2_51 100 105 2.16e-15
C2_52 103 105 2.16e-15
R2_6 101 100 0.001
C2_61 101 105 8.4e-16
C2_62 100 105 8.4e-16
R2_7 102 101 0.001
C2_71 102 105 2.4e-16
C2_72 101 105 2.4e-16
R2_8 99 102 0.001
C2_81 99 105 3.6e-16
C2_82 102 105 3.6e-16
R2_9 97 99 0.1
C2_91 97 105 2.16e-15
C2_92 99 105 2.16e-15
R2_10 95 97 0.001
C2_101 95 105 8.4e-16
C2_102 97 105 8.4e-16
R2_11 96 95 0.001
C2_111 96 105 2.4e-16
C2_112 95 105 2.4e-16
R2_12 94 96 0.001
C2_121 94 105 3.6e-16
C2_122 96 105 3.6e-16
R2_13 94 105 0.001
C2_131 94 105 1.2e-15
C2_132 105 105 1.2e-15
R2_14 91 105 0.001
C2_141 91 105 9.6e-16
C2_142 105 105 9.6e-16
R2_15 92 91 0.001
C2_151 92 105 1.08e-15
C2_152 91 105 1.08e-15
R1_1 108 109 0.001
R1_2 119 120 0.001
R1_3 128 127 0.001
R1_4 122 121 0.001
R1_5 128 129 0.001
R1_6 124 123 0.001
R1_7 136 135 0.001
R1_8 131 130 0.001
R1_9 116 115 0.001
R1_10 135 137 0.001
R1_11 131 132 0.001
R1_12 134 133 0.001
R1_13 151 152 0.001
R1_14 145 146 0.001
R1_15 139 138 0.001
R1_16 117 118 0.001
R1_17 138 140 0.001
R1_18 144 143 0.001
R1_19 149 150 0.001
R1_20 148 147 0.001
R1_21 148 153 500
C1_211 148 105 1.575e-15
C1_212 153 105 1.575e-15
R1_22 141 148 550
C1_221 141 105 1.65e-15
C1_222 148 105 1.65e-15
R1_23 149 154 500
C1_231 149 105 1.575e-15
C1_232 154 105 1.575e-15
R1_24 142 149 550
C1_241 142 105 1.65e-15
C1_242 149 105 1.65e-15
R1_25 147 156 0.6
C1_251 147 105 1.75e-15
C1_252 156 105 1.75e-15
R1_26 140 147 0.9
C1_261 140 105 2.52e-15
C1_262 147 105 2.52e-15
R1_27 150 157 0.6
C1_271 150 105 1.75e-15
C1_272 157 105 1.75e-15
R1_28 143 150 0.9
C1_281 143 105 2.52e-15
C1_282 150 105 2.52e-15
R1_29 117 126 550
C1_291 117 105 1.65e-15
C1_292 126 105 1.65e-15
R1_30 113 117 500
C1_301 113 105 1.575e-15
C1_302 117 105 1.575e-15
R1_31 138 144 0.35
C1_311 138 105 1.8e-15
C1_312 144 105 1.8e-15
R1_32 118 133 0.9
C1_321 118 105 2.52e-15
C1_322 133 105 2.52e-15
R1_33 114 118 0.6
C1_331 114 105 1.75e-15
C1_332 118 105 1.75e-15
R1_34 132 139 0.5
C1_341 132 105 2.4e-15
C1_342 139 105 2.4e-15
R1_35 152 155 0.001
C1_351 152 105 2.1e-16
C1_352 155 105 2.1e-16
R1_36 146 152 1
C1_361 146 105 2.8e-15
C1_362 152 105 2.8e-15
R1_37 137 146 0.4
C1_371 137 105 1.26e-15
C1_372 146 105 1.26e-15
R1_38 116 125 550
C1_381 116 105 1.65e-15
C1_382 125 105 1.65e-15
R1_39 112 116 500
C1_391 112 105 1.575e-15
C1_392 116 105 1.575e-15
R1_40 131 134 0.35
C1_401 131 105 1.8e-15
C1_402 134 105 1.8e-15
R1_41 123 130 0.2
C1_411 123 105 7e-16
C1_412 130 105 7e-16
R1_42 115 123 0.6
C1_421 115 105 1.82e-15
C1_422 123 105 1.82e-15
R1_43 111 115 0.6
C1_431 111 105 1.75e-15
C1_432 115 105 1.75e-15
R1_44 129 136 0.5
C1_441 129 105 2.4e-15
C1_442 136 105 2.4e-15
R1_45 122 124 0.25
C1_451 122 105 1.2e-15
C1_452 124 105 1.2e-15
R1_46 121 127 0.2
C1_461 121 105 7e-16
C1_462 127 105 7e-16
R1_47 120 121 0.2
C1_471 120 105 5.6e-16
C1_472 121 105 5.6e-16
R1_48 109 120 1
C1_481 109 105 2.8e-15
C1_482 120 105 2.8e-15
R1_49 110 109 0.001
C1_491 110 105 2.1e-16
C1_492 109 105 2.1e-16
.ends fo4_eq2

