
.include nand2_teste4.spi

* INTERF a b vdd vss y

X1 10 11 40 30 20 nand2_teste4

V1 10 30 dc 0.0V
V2 11 30 dc 1.8V
Vdd 40 30 1.8V
Vss 30 0 0.0V

.model tp pmos level = 54
.model tn nmos level = 54

.dc V1 0 1.8 0.001
.end

