* Spice description of mux2
* Spice driver version -1218375111
* Date ( dd/mm/yyyy hh:mm:ss ):  5/11/2020 at 15:51:34

* INTERF a0 a1 n_s s vdd vss y 


.subckt mux2 63 72 44 25 3 51 80 
* NET 3 = vdd
* NET 25 = s
* NET 44 = n_s
* NET 51 = vss
* NET 63 = a0
* NET 72 = a1
* NET 80 = y
Mtr_00004 64 21 82 3 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 71 40 84 3 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 60 31 76 51 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 68 13 79 51 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R7_1 5 4 0.001
R7_2 1 3 0.001
R7_3 3 6 0.001
C7_31 3 51 8.4e-16
C7_32 6 51 8.4e-16
R7_4 2 3 0.1
C7_41 2 51 2.76e-15
C7_42 3 51 2.76e-15
R7_5 4 8 0.1
C7_51 4 51 2.76e-15
C7_52 8 51 2.76e-15
R7_6 7 4 0.001
C7_61 7 51 8.4e-16
C7_62 4 51 8.4e-16
R7_7 6 7 0.001
C7_71 6 51 2.4e-16
C7_72 7 51 2.4e-16
R6_1 19 14 0.001
R6_2 14 15 0.001
R6_3 15 16 0.001
R6_4 12 11 0.001
R6_5 23 22 0.001
R6_6 22 24 0.001
R6_7 27 26 0.001
R6_8 21 27 300
C6_81 21 51 9.75e-16
C6_82 27 51 9.75e-16
R6_9 26 28 0.2
C6_91 26 51 2.875e-16
C6_92 28 51 2.875e-16
R6_10 25 26 0.3
C6_101 25 51 3.45e-16
C6_102 26 51 3.45e-16
R6_11 24 25 0.5
C6_111 24 51 5.75e-16
C6_112 25 51 5.75e-16
R6_12 12 23 0.35
C6_121 12 51 1.8e-15
C6_122 23 51 1.8e-15
R6_13 11 15 0.35
C6_131 11 51 1.68e-15
C6_132 15 51 1.68e-15
R6_14 17 13 200
C6_141 17 51 6e-16
C6_142 13 51 6e-16
R6_15 14 20 0.5
C6_151 14 51 5.75e-16
C6_152 20 51 5.75e-16
R6_16 18 14 0.6
C6_161 18 51 6.9e-16
C6_162 14 51 6.9e-16
R6_17 13 19 200
C6_171 13 51 6.75e-16
C6_172 19 51 6.75e-16
R5_1 35 34 0.001
R5_2 37 36 0.001
R5_3 39 38 0.001
R5_4 42 41 0.001
R5_5 41 43 0.001
R5_6 46 45 0.001
R5_7 40 46 300
C5_71 40 51 9.75e-16
C5_72 46 51 9.75e-16
R5_8 45 47 0.2
C5_81 45 51 2.875e-16
C5_82 47 51 2.875e-16
R5_9 44 45 0.3
C5_91 44 51 3.45e-16
C5_92 45 51 3.45e-16
R5_10 43 44 0.5
C5_101 43 51 5.75e-16
C5_102 44 51 5.75e-16
R5_11 39 42 0.25
C5_111 39 51 1.2e-15
C5_112 42 51 1.2e-15
R5_12 37 38 0.35
C5_121 37 51 1.68e-15
C5_122 38 51 1.68e-15
R5_13 34 36 0.4
C5_131 34 51 4.6e-16
C5_132 36 51 4.6e-16
R5_14 32 34 0.6
C5_141 32 51 7.475e-16
C5_142 34 51 7.475e-16
R5_15 31 35 200
C5_151 31 51 6.75e-16
C5_152 35 51 6.75e-16
R5_16 33 31 200
C5_161 33 51 6e-16
C5_162 31 51 6e-16
R4_1 57 52 0.001
R4_2 56 51 0.001
R4_3 51 53 0.001
C4_31 51 51 8.4e-16
C4_32 53 51 8.4e-16
R4_4 50 51 0.1
C4_41 50 51 2.76e-15
C4_42 51 51 2.76e-15
R4_5 52 55 0.1
C4_51 52 51 2.76e-15
C4_52 55 51 2.76e-15
R4_6 54 52 0.001
C4_61 54 51 8.4e-16
C4_62 52 51 8.4e-16
R4_7 53 54 0.001
C4_71 53 51 2.4e-16
C4_72 54 51 2.4e-16
R3_1 60 61 0.001
R3_2 64 63 0.001
R3_3 63 65 0.4
C3_31 63 51 1.365e-15
C3_32 65 51 1.365e-15
R3_4 61 63 0.9
C3_41 61 51 2.765e-15
C3_42 63 51 2.765e-15
R3_5 62 61 0.001
C3_51 62 51 2.1e-16
C3_52 61 51 2.1e-16
R2_1 68 69 0.001
R2_2 71 72 0.001
R2_3 72 73 0.4
C2_31 72 51 1.365e-15
C2_32 73 51 1.365e-15
R2_4 69 72 0.9
C2_41 69 51 2.765e-15
C2_42 72 51 2.765e-15
R2_5 70 69 0.001
C2_51 70 51 2.1e-16
C2_52 69 51 2.1e-16
R1_1 79 80 0.001
R1_2 80 81 0.001
R1_3 84 85 0.001
R1_4 78 77 0.001
R1_5 77 76 0.001
R1_6 82 83 0.001
R1_7 83 86 0.1
C1_71 83 51 1.725e-16
C1_72 86 51 1.725e-16
R1_8 77 83 2
C1_81 77 51 2.3575e-15
C1_82 83 51 2.3575e-15
R1_9 78 81 0.1
C1_91 78 51 4.8e-16
C1_92 81 51 4.8e-16
R1_10 85 87 0.1
C1_101 85 51 1.725e-16
C1_102 87 51 1.725e-16
R1_11 80 85 2
C1_111 80 51 2.3575e-15
C1_112 85 51 2.3575e-15
.ends mux2

