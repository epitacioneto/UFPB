* Spice description of nand2_teste2
* Spice driver version -1218080199
* Date ( dd/mm/yyyy hh:mm:ss ):  3/11/2020 at 18:12:01

* INTERF a b vdd vss y 


.subckt nand2_teste2 1 11 21 39 33 
* NET 1 = a
* NET 11 = b
* NET 21 = vdd
* NET 33 = y
* NET 39 = vss
Mtr_00004 34 12 20 21 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00003 34 7 19 21 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00002 28 5 40 39 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 28 10 31 39 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
R5_1 3 2 0.001
R5_2 2 6 0.9
C5_21 2 39 2.59e-15
C5_22 6 39 2.59e-15
R5_3 1 2 0.1
C5_31 1 39 2.8e-16
C5_32 2 39 2.8e-16
R5_4 4 1 0.5
C5_41 4 39 1.47e-15
C5_42 1 39 1.47e-15
R5_5 3 7 450
C5_51 3 39 1.35e-15
C5_52 7 39 1.35e-15
R5_6 5 3 500
C5_61 5 39 1.575e-15
C5_62 3 39 1.575e-15
R4_1 15 14 0.001
R4_2 14 16 0.9
C4_21 14 39 2.59e-15
C4_22 16 39 2.59e-15
R4_3 11 14 0.1
C4_31 11 39 2.8e-16
C4_32 14 39 2.8e-16
R4_4 13 12 450
C4_41 13 39 1.35e-15
C4_42 12 39 1.35e-15
R4_5 10 13 450
C4_51 10 39 1.425e-15
C4_52 13 39 1.425e-15
R4_6 13 15 200
C4_61 13 39 6e-16
C4_62 15 39 6e-16
R3_1 19 21 0.001
R3_2 20 24 0.001
R3_3 24 25 0.001
C3_31 24 39 1.08e-15
C3_32 25 39 1.08e-15
R3_4 23 24 0.1
C3_41 23 39 1.44e-15
C3_42 24 39 1.44e-15
R3_5 21 23 0.1
C3_51 21 39 1.44e-15
C3_52 23 39 1.44e-15
R3_6 22 21 0.001
C3_61 22 39 1.08e-15
C3_62 21 39 1.08e-15
R2_1 31 32 0.001
R2_2 28 29 0.001
R2_3 34 35 0.001
R2_4 35 36 0.2
C2_41 35 39 6.3e-16
C2_42 36 39 6.3e-16
R2_5 33 35 0.8
C2_51 33 39 2.24e-15
C2_52 35 39 2.24e-15
R2_6 29 33 0.4
C2_61 29 39 1.26e-15
C2_62 33 39 1.26e-15
R2_7 30 29 0.001
C2_71 30 39 2.1e-16
C2_72 29 39 2.1e-16
R2_8 29 32 0.6
C2_81 29 39 6.9e-16
C2_82 32 39 6.9e-16
R1_1 40 39 0.001
R1_2 41 39 0.001
C1_21 41 39 1.08e-15
C1_22 39 39 1.08e-15
R1_3 43 44 0.001
C1_31 43 39 1.2e-15
C1_32 44 39 1.2e-15
R1_4 42 43 0.001
C1_41 42 39 1.32e-15
C1_42 43 39 1.32e-15
R1_5 39 42 0.1
C1_51 39 39 1.44e-15
C1_52 42 39 1.44e-15
.ends nand2_teste2

