* Spice description of nand2_teste3
* Spice driver version -1218018759
* Date ( dd/mm/yyyy hh:mm:ss ):  3/11/2020 at 18:53:56

* INTERF a b vdd vss y 


.subckt nand2_teste3 10 2 21 31 43 
* NET 2 = b
* NET 10 = a
* NET 21 = vdd
* NET 31 = vss
* NET 43 = y
Mtr_00004 44 16 19 21 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 44 3 20 21 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 28 14 32 31 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 28 1 40 31 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R6_1 6 5 0.001
R6_2 4 3 450
C6_21 4 31 1.425e-15
C6_22 3 31 1.425e-15
R6_3 1 4 500
C6_31 1 31 1.575e-15
C6_32 4 31 1.575e-15
R6_4 5 7 0.9
C6_41 5 31 2.59e-15
C6_42 7 31 2.59e-15
R6_5 2 5 0.1
C6_51 2 31 2.8e-16
C6_52 5 31 2.8e-16
R6_6 4 6 150
C6_61 4 31 4.5e-16
C6_62 6 31 4.5e-16
R5_1 12 11 0.001
R5_2 11 15 0.9
C5_21 11 31 2.59e-15
C5_22 15 31 2.59e-15
R5_3 10 11 0.1
C5_31 10 31 2.8e-16
C5_32 11 31 2.8e-16
R5_4 13 10 0.5
C5_41 13 31 1.47e-15
C5_42 10 31 1.47e-15
R5_5 12 16 450
C5_51 12 31 1.425e-15
C5_52 16 31 1.425e-15
R5_6 14 12 500
C5_61 14 31 1.575e-15
C5_62 12 31 1.575e-15
R4_1 20 24 0.001
R4_2 19 21 0.001
R4_3 24 25 0.001
C4_31 24 31 1.32e-15
C4_32 25 31 1.32e-15
R4_4 23 24 0.001
C4_41 23 31 1.2e-15
C4_42 24 31 1.2e-15
R4_5 21 23 0.1
C4_51 21 31 1.44e-15
C4_52 23 31 1.44e-15
R4_6 22 21 0.001
C4_61 22 31 1.08e-15
C4_62 21 31 1.08e-15
R2_1 32 31 0.001
R2_2 33 31 0.001
C2_21 33 31 1.08e-15
C2_22 31 31 1.08e-15
R2_3 35 36 0.001
C2_31 35 31 1.2e-15
C2_32 36 31 1.2e-15
R2_4 34 35 0.001
C2_41 34 31 1.08e-15
C2_42 35 31 1.08e-15
R2_5 31 34 0.1
C2_51 31 31 1.68e-15
C2_52 34 31 1.68e-15
R1_1 40 41 0.001
R1_2 44 45 0.001
R1_3 45 46 0.4
C1_31 45 31 1.33e-15
C1_32 46 31 1.33e-15
R1_4 43 45 0.5
C1_41 43 31 1.54e-15
C1_42 45 31 1.54e-15
R1_5 39 43 0.5
C1_51 39 31 1.4e-15
C1_52 43 31 1.4e-15
R1_6 41 42 0.1
C1_61 41 31 1.725e-16
C1_62 42 31 1.725e-16
R1_7 39 41 0.5
C1_71 39 31 5.75e-16
C1_72 41 31 5.75e-16
.ends nand2_teste3

