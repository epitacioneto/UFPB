* Spice description of fo4+gordo
* Spice driver version -1217572295
* Date ( dd/mm/yyyy hh:mm:ss ): 19/10/2020 at 15:09:11

* INTERF a vdd vss vss1 y 


.subckt fo4+gordo 42 61 123 5 90 
* NET 5 = vss1
* NET 42 = a
* NET 61 = vdd
* NET 90 = y
* NET 123 = vss
Mtr_00010 14 97 63 61 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 33 77 48 61 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 22 96 62 61 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 129 74 47 61 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 79 43 46 61 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00005 17 104 2 123 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00004 30 71 116 123 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 25 102 1 123 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 126 69 111 123 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 66 41 108 123 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
R9_1 1 3 0.001
R9_2 2 8 0.001
R9_3 10 11 0.001
C9_31 10 123 6e-16
C9_32 11 123 6e-16
R9_4 8 10 0.1
C9_41 8 123 2.16e-15
C9_42 10 123 2.16e-15
R9_5 9 8 0.001
C9_51 9 123 8.4e-16
C9_52 8 123 8.4e-16
R9_6 7 9 0.001
C9_61 7 123 2.4e-16
C9_62 9 123 2.4e-16
R9_7 6 7 0.001
C9_71 6 123 3.6e-16
C9_72 7 123 3.6e-16
R9_8 6 5 0.001
C9_81 6 123 1.2e-15
C9_82 5 123 1.2e-15
R9_9 3 5 0.001
C9_91 3 123 9.6e-16
C9_92 5 123 9.6e-16
R9_10 4 3 0.001
C9_101 4 123 1.08e-15
C9_102 3 123 1.08e-15
R8_1 17 18 0.001
R8_2 14 15 0.001
R8_3 18 19 0.001
C8_31 18 123 2.1e-16
C8_32 19 123 2.1e-16
R8_4 15 18 1
C8_41 15 123 2.8e-15
C8_42 18 123 2.8e-15
R8_5 16 15 0.4
C8_51 16 123 1.33e-15
C8_52 15 123 1.33e-15
R7_1 25 26 0.001
R7_2 22 23 0.001
R7_3 26 27 0.001
C7_31 26 123 2.1e-16
C7_32 27 123 2.1e-16
R7_4 23 26 1
C7_41 23 123 2.8e-15
C7_42 26 123 2.8e-15
R7_5 24 23 0.4
C7_51 24 123 1.33e-15
C7_52 23 123 1.33e-15
R6_1 30 31 0.001
R6_2 33 34 0.001
R6_3 34 35 0.4
C6_31 34 123 1.33e-15
C6_32 35 123 1.33e-15
R6_4 31 34 1
C6_41 31 123 2.8e-15
C6_42 34 123 2.8e-15
R6_5 32 31 0.001
C6_51 32 123 2.1e-16
C6_52 31 123 2.1e-16
R5_1 39 38 0.001
R5_2 38 42 0.9
C5_21 38 123 2.52e-15
C5_22 42 123 2.52e-15
R5_3 40 38 0.6
C5_31 40 123 1.75e-15
C5_32 38 123 1.75e-15
R5_4 39 43 650
C5_41 39 123 2.025e-15
C5_42 43 123 2.025e-15
R5_5 41 39 550
C5_51 41 123 1.725e-15
C5_52 39 123 1.725e-15
R4_1 46 49 0.001
R4_2 47 52 0.001
R4_3 62 52 0.001
R4_4 48 58 0.001
R4_5 63 58 0.001
R4_6 59 60 0.001
C4_61 59 123 2.145e-15
C4_62 60 123 2.145e-15
R4_7 58 59 0.001
C4_71 58 123 2.34e-15
C4_72 59 123 2.34e-15
R4_8 56 58 0.001
C4_81 56 123 1.365e-15
C4_82 58 123 1.365e-15
R4_9 57 56 0.001
C4_91 57 123 3.9e-16
C4_92 56 123 3.9e-16
R4_10 55 57 0.001
C4_101 55 123 1.755e-15
C4_102 57 123 1.755e-15
R4_11 52 55 0.001
C4_111 52 123 2.34e-15
C4_112 55 123 2.34e-15
R4_12 53 52 0.001
C4_121 53 123 1.365e-15
C4_122 52 123 1.365e-15
R4_13 54 53 0.001
C4_131 54 123 3.9e-16
C4_132 53 123 3.9e-16
R4_14 51 54 0.001
C4_141 51 123 1.08e-15
C4_142 54 123 1.08e-15
R4_15 51 61 0.001
C4_151 51 123 7.2e-16
C4_152 61 123 7.2e-16
R4_16 49 61 0.001
C4_161 49 123 7.2e-16
C4_162 61 123 7.2e-16
R4_17 50 49 0.001
C4_171 50 123 1.08e-15
C4_172 49 123 1.08e-15
R3_1 66 67 0.001
R3_2 79 80 0.001
R3_3 82 81 0.001
R3_4 84 83 0.001
R3_5 86 85 0.001
R3_6 73 75 0.001
R3_7 86 87 0.001
R3_8 89 88 0.001
R3_9 92 91 0.001
R3_10 76 78 0.001
R3_11 91 93 0.001
R3_12 95 94 0.001
R3_13 100 101 0.001
R3_14 98 99 0.001
R3_15 98 102 500
C3_151 98 123 1.575e-15
C3_152 102 123 1.575e-15
R3_16 96 98 550
C3_161 96 123 1.65e-15
C3_162 98 123 1.65e-15
R3_17 100 104 500
C3_171 100 123 1.575e-15
C3_172 104 123 1.575e-15
R3_18 97 100 550
C3_181 97 123 1.65e-15
C3_182 100 123 1.65e-15
R3_19 99 103 0.6
C3_191 99 123 1.75e-15
C3_192 103 123 1.75e-15
R3_20 93 99 0.9
C3_201 93 123 2.52e-15
C3_202 99 123 2.52e-15
R3_21 101 105 0.6
C3_211 101 123 1.75e-15
C3_212 105 123 1.75e-15
R3_22 94 101 0.9
C3_221 94 123 2.52e-15
C3_222 101 123 2.52e-15
R3_23 76 77 550
C3_231 76 123 1.65e-15
C3_232 77 123 1.65e-15
R3_24 71 76 500
C3_241 71 123 1.575e-15
C3_242 76 123 1.575e-15
R3_25 91 95 0.35
C3_251 91 123 1.8e-15
C3_252 95 123 1.8e-15
R3_26 78 88 0.9
C3_261 78 123 2.52e-15
C3_262 88 123 2.52e-15
R3_27 72 78 0.6
C3_271 72 123 1.75e-15
C3_272 78 123 1.75e-15
R3_28 87 92 0.5
C3_281 87 123 2.4e-15
C3_282 92 123 2.4e-15
R3_29 73 74 550
C3_291 73 123 1.65e-15
C3_292 74 123 1.65e-15
R3_30 69 73 500
C3_301 69 123 1.575e-15
C3_302 73 123 1.575e-15
R3_31 86 89 0.35
C3_311 86 123 1.8e-15
C3_312 89 123 1.8e-15
R3_32 83 85 0.2
C3_321 83 123 7e-16
C3_322 85 123 7e-16
R3_33 75 83 0.6
C3_331 75 123 1.82e-15
C3_332 83 123 1.82e-15
R3_34 70 75 0.6
C3_341 70 123 1.75e-15
C3_342 75 123 1.75e-15
R3_35 82 84 0.25
C3_351 82 123 1.2e-15
C3_352 84 123 1.2e-15
R3_36 81 90 0.2
C3_361 81 123 7e-16
C3_362 90 123 7e-16
R3_37 80 81 0.2
C3_371 80 123 5.6e-16
C3_372 81 123 5.6e-16
R3_38 67 80 1
C3_381 67 123 2.8e-15
C3_382 80 123 2.8e-15
R3_39 68 67 0.001
C3_391 68 123 2.1e-16
C3_392 67 123 2.1e-16
R2_1 111 115 0.001
R2_2 116 118 0.001
R2_3 108 109 0.001
R2_4 112 113 0.001
C2_41 112 123 3.6e-16
C2_42 113 123 3.6e-16
R2_5 112 123 0.001
C2_51 112 123 1.2e-15
C2_52 123 123 1.2e-15
R2_6 109 123 0.001
C2_61 109 123 9.6e-16
C2_62 123 123 9.6e-16
R2_7 110 109 0.001
C2_71 110 123 1.08e-15
C2_72 109 123 1.08e-15
R2_8 121 122 0.001
C2_81 121 123 6e-16
C2_82 122 123 6e-16
R2_9 118 121 0.1
C2_91 118 123 2.16e-15
C2_92 121 123 2.16e-15
R2_10 119 118 0.001
C2_101 119 123 8.4e-16
C2_102 118 123 8.4e-16
R2_11 120 119 0.001
C2_111 120 123 2.4e-16
C2_112 119 123 2.4e-16
R2_12 117 120 0.001
C2_121 117 123 3.6e-16
C2_122 120 123 3.6e-16
R2_13 115 117 0.1
C2_131 115 123 2.16e-15
C2_132 117 123 2.16e-15
R2_14 114 115 0.001
C2_141 114 123 8.4e-16
C2_142 115 123 8.4e-16
R2_15 113 114 0.001
C2_151 113 123 2.4e-16
C2_152 114 123 2.4e-16
R1_1 126 127 0.001
R1_2 129 130 0.001
R1_3 130 131 0.4
C1_31 130 123 1.33e-15
C1_32 131 123 1.33e-15
R1_4 127 130 1
C1_41 127 123 2.8e-15
C1_42 130 123 2.8e-15
R1_5 128 127 0.001
C1_51 128 123 2.1e-16
C1_52 127 123 2.1e-16
.ends fo4+gordo

