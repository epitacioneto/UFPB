* Spice description of latch_d_roteado
* Spice driver version -1218387399
* Date ( dd/mm/yyyy hh:mm:ss ): 19/11/2020 at 15:23:45

* INTERF a ck q vdd vss 


.subckt latch_d_roteado 7 8 5 12 3 
* NET 3 = vss
* NET 4 = q_b
* NET 5 = q
* NET 6 = b
* NET 7 = a
* NET 8 = ck
* NET 12 = vdd
Mtr_00016 12 11 5 12 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00015 13 7 12 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 9 8 12 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 10 8 11 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00012 11 9 13 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 12 6 10 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 4 5 12 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 6 4 12 12 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 3 7 2 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 2 8 11 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 3 8 9 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 11 9 1 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 1 6 3 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 5 11 3 3 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 3 5 4 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 3 4 6 3 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C11 3 3 1.0176e-13
C10 4 3 4.897e-14
C9 5 3 5.101e-14
C8 6 3 6.088e-14
C7 7 3 3.309e-14
C6 8 3 4.268e-14
C5 9 3 2.356e-14
C3 11 3 1.932e-14
C2 12 3 1.1044e-13
.ends latch_d_roteado

