* Spice description of tristate
* Spice driver version -1217535431
* Date ( dd/mm/yyyy hh:mm:ss ):  5/11/2020 at 15:10:37

* INTERF a enable n_enable vdd vss y 


.subckt tristate 28 15 8 2 20 39 
* NET 2 = vdd
* NET 8 = n_enable
* NET 15 = enable
* NET 20 = vss
* NET 28 = a
* NET 39 = y
Mtr_00002 29 7 37 2 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 25 13 34 20 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R6_1 3 2 0.001
R6_2 2 4 0.001
C6_21 2 20 1.08e-15
C6_22 4 20 1.08e-15
R6_3 1 2 0.1
C6_31 1 20 2.76e-15
C6_32 2 20 2.76e-15
R5_1 9 8 0.001
R5_2 10 9 150
C5_21 10 20 4.5e-16
C5_22 9 20 4.5e-16
R5_3 7 10 300
C5_31 7 20 9.75e-16
C5_32 10 20 9.75e-16
R4_1 16 15 0.001
R4_2 14 13 200
C4_21 14 20 6e-16
C4_22 13 20 6e-16
R4_3 13 16 200
C4_31 13 20 6.75e-16
C4_32 16 20 6.75e-16
R3_1 21 20 0.001
R3_2 20 22 0.001
C3_21 20 20 1.08e-15
C3_22 22 20 1.08e-15
R3_3 19 20 0.1
C3_31 19 20 2.76e-15
C3_32 20 20 2.76e-15
R2_1 25 26 0.001
R2_2 29 30 0.001
R2_3 30 31 0.4
C2_31 30 20 1.33e-15
C2_32 31 20 1.33e-15
R2_4 28 30 0.1
C2_41 28 20 4.2e-16
C2_42 30 20 4.2e-16
R2_5 26 28 0.8
C2_51 26 20 2.38e-15
C2_52 28 20 2.38e-15
R2_6 27 26 0.001
C2_61 27 20 2.1e-16
C2_62 26 20 2.1e-16
R1_1 34 35 0.001
R1_2 37 38 0.001
R1_3 38 40 0.1
C1_31 38 20 1.725e-16
C1_32 40 20 1.725e-16
R1_4 39 38 0.3
C1_41 39 20 3.45e-16
C1_42 38 20 3.45e-16
R1_5 35 39 1.7
C1_51 35 20 1.955e-15
C1_52 39 20 1.955e-15
R1_6 36 35 0.1
C1_61 36 20 1.725e-16
C1_62 35 20 1.725e-16
.ends tristate

