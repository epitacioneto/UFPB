
.include fo4_inveq_s.spi
.include inversor_equilibrado.spi

* a vdd vss y 
X1 20 10 30 40 fo4_inveq_s
X2 20 10 30 41 inversor_equilibrado

V1 10 30 1.8V DC
V2 30 0 0V DC
V3 20 30 pulse(0V 1.8V 2ns 1ps 1ps 2ns 4ns)

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.001ns 8ns

.end
