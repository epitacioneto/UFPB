* Spice description of tran_passagem
* Spice driver version -1217768903
* Date ( dd/mm/yyyy hh:mm:ss ):  3/11/2020 at 14:35:10

* INTERF a enable vdd vss y1 y2 


.subckt tran_passagem 59 9 14 41 24 53 
* NET 9 = enable
* NET 14 = vdd
* NET 24 = y1
* NET 41 = vss
* NET 53 = y2
* NET 59 = a
Mtr_00004 60 34 23 14 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 32 6 13 14 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 56 4 51 41 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 29 1 42 41 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R7_1 8 7 0.001
R7_2 9 10 0.2
C7_21 9 41 7.7e-16
C7_22 10 41 7.7e-16
R7_3 7 9 0.6
C7_31 7 41 1.82e-15
C7_32 9 41 1.82e-15
R7_4 2 7 0.6
C7_41 2 41 1.75e-15
C7_42 7 41 1.75e-15
R7_5 8 6 450
C7_51 8 41 1.425e-15
C7_52 6 41 1.425e-15
R7_6 1 8 500
C7_61 1 41 1.575e-15
C7_62 8 41 1.575e-15
R7_7 3 1 150
C7_71 3 41 5.25e-16
C7_72 1 41 5.25e-16
R7_8 3 5 800
C7_81 3 41 2.4e-15
C7_82 5 41 2.4e-15
R7_9 5 4 150
C7_91 5 41 5.25e-16
C7_92 4 41 5.25e-16
R6_1 13 14 0.001
R6_2 19 18 0.001
R6_3 18 20 0.001
C6_31 18 41 1.08e-15
C6_32 20 41 1.08e-15
R6_4 16 18 0.1
C6_41 16 41 2.52e-15
C6_42 18 41 2.52e-15
R6_5 17 16 0.001
C6_51 17 41 2.4e-16
C6_52 16 41 2.4e-16
R6_6 14 17 0.1
C6_61 14 41 2.52e-15
C6_62 17 41 2.52e-15
R6_7 15 14 0.001
C6_71 15 41 1.08e-15
C6_72 14 41 1.08e-15
R5_1 23 25 0.001
R5_2 25 26 0.1
C5_21 25 41 1.725e-16
C5_22 26 41 1.725e-16
R5_3 24 25 0.3
C5_31 24 41 3.45e-16
C5_32 25 41 3.45e-16
R4_1 29 30 0.001
R4_2 36 35 0.001
R4_3 32 33 0.001
R4_4 34 37 300
C4_41 34 41 9.75e-16
C4_42 37 41 9.75e-16
R4_5 36 37 650
C4_51 36 41 1.95e-15
C4_52 37 41 1.95e-15
R4_6 35 38 0.1
C4_61 35 41 3.5e-16
C4_62 38 41 3.5e-16
R4_7 33 35 0.3
C4_71 33 41 9.8e-16
C4_72 35 41 9.8e-16
R4_8 30 33 1
C4_81 30 41 2.8e-15
C4_82 33 41 2.8e-15
R4_9 31 30 0.001
C4_91 31 41 2.1e-16
C4_92 30 41 2.1e-16
R3_1 42 41 0.001
R3_2 47 46 0.001
R3_3 46 48 0.001
C3_31 46 41 1.08e-15
C3_32 48 41 1.08e-15
R3_4 44 46 0.1
C3_41 44 41 2.52e-15
C3_42 46 41 2.52e-15
R3_5 45 44 0.001
C3_51 45 41 2.4e-16
C3_52 44 41 2.4e-16
R3_6 41 45 0.1
C3_61 41 41 2.52e-15
C3_62 45 41 2.52e-15
R3_7 43 41 0.001
C3_71 43 41 1.08e-15
C3_72 41 41 1.08e-15
R2_1 51 52 0.001
R2_2 52 53 0.3
C2_21 52 41 3.45e-16
C2_22 53 41 3.45e-16
R1_1 56 57 0.001
R1_2 60 61 0.001
R1_3 61 62 0.4
C1_31 61 41 1.33e-15
C1_32 62 41 1.33e-15
R1_4 59 61 0.3
C1_41 59 41 8.4e-16
C1_42 61 41 8.4e-16
R1_5 57 59 0.7
C1_51 57 41 1.96e-15
C1_52 59 41 1.96e-15
R1_6 58 57 0.001
C1_61 58 41 2.1e-16
C1_62 57 41 2.1e-16
.ends tran_passagem

