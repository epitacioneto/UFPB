
.include nand2_teste4.spi

* INTERF a b vdd vss y

X1 10 11 40 30 20 nand2_teste4

V1 10 30 pulse(0 1.8V 3ns 1ps 1ps 4ns 8ns)
V2 11 30 pulse(0 1.8V 1ns 1ps 1ps 2ns 5ns)
Vdd 40 30 1.8V
Vss 30 0 0.0V

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.001ns 20ns
.end

