* Spice description of fo4_gordo2
* Spice driver version -1217781191
* Date ( dd/mm/yyyy hh:mm:ss ): 19/10/2020 at 22:36:03

* INTERF a vdd vss vss1 y 


.subckt fo4_gordo2 47 77 149 16 101 
* NET 16 = vss1
* NET 47 = a
* NET 77 = vdd
* NET 101 = y
* NET 149 = vss
Mtr_00012 109 51 76 77 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00011 19 120 79 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 38 100 63 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 27 119 78 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 155 99 62 77 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 93 50 61 77 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 125 58 1 149 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00005 22 128 3 149 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00004 35 87 142 149 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 30 127 2 149 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 152 86 137 149 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 82 46 134 149 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
R9_1 1 4 0.001
R9_2 2 9 0.001
R9_3 3 11 0.001
R9_4 14 15 0.001
C9_41 14 149 6e-16
C9_42 15 149 6e-16
R9_5 11 14 0.1
C9_51 11 149 2.16e-15
C9_52 14 149 2.16e-15
R9_6 12 11 0.001
C9_61 12 149 8.4e-16
C9_62 11 149 8.4e-16
R9_7 13 12 0.001
C9_71 13 149 2.4e-16
C9_72 12 149 2.4e-16
R9_8 10 13 0.001
C9_81 10 149 3.6e-16
C9_82 13 149 3.6e-16
R9_9 10 16 0.001
C9_91 10 149 1.2e-15
C9_92 16 149 1.2e-15
R9_10 9 16 0.001
C9_101 9 149 9.6e-16
C9_102 16 149 9.6e-16
R9_11 7 9 0.001
C9_111 7 149 8.4e-16
C9_112 9 149 8.4e-16
R9_12 8 7 0.001
C9_121 8 149 2.4e-16
C9_122 7 149 2.4e-16
R9_13 6 8 0.001
C9_131 6 149 3.6e-16
C9_132 8 149 3.6e-16
R9_14 4 6 0.1
C9_141 4 149 2.16e-15
C9_142 6 149 2.16e-15
R9_15 5 4 0.001
C9_151 5 149 1.08e-15
C9_152 4 149 1.08e-15
R8_1 22 23 0.001
R8_2 19 20 0.001
R8_3 23 24 0.001
C8_31 23 149 2.1e-16
C8_32 24 149 2.1e-16
R8_4 20 23 1
C8_41 20 149 2.8e-15
C8_42 23 149 2.8e-15
R8_5 21 20 0.4
C8_51 21 149 1.33e-15
C8_52 20 149 1.33e-15
R7_1 30 31 0.001
R7_2 27 28 0.001
R7_3 31 32 0.001
C7_31 31 149 2.1e-16
C7_32 32 149 2.1e-16
R7_4 28 31 1
C7_41 28 149 2.8e-15
C7_42 31 149 2.8e-15
R7_5 29 28 0.4
C7_51 29 149 1.33e-15
C7_52 28 149 1.33e-15
R6_1 35 36 0.001
R6_2 38 39 0.001
R6_3 39 40 0.4
C6_31 39 149 1.33e-15
C6_32 40 149 1.33e-15
R6_4 36 39 1
C6_41 36 149 2.8e-15
C6_42 39 149 2.8e-15
R6_5 37 36 0.001
C6_51 37 149 2.1e-16
C6_52 36 149 2.1e-16
R5_1 44 43 0.001
R5_2 48 47 0.001
R5_3 48 49 0.001
R5_4 53 52 0.001
R5_5 52 54 0.001
R5_6 56 55 0.001
R5_7 56 58 550
C5_71 56 149 1.725e-15
C5_72 58 149 1.725e-15
R5_8 51 56 650
C5_81 51 149 2.025e-15
C5_82 56 149 2.025e-15
R5_9 55 57 0.6
C5_91 55 149 1.75e-15
C5_92 57 149 1.75e-15
R5_10 54 55 0.9
C5_101 54 149 2.52e-15
C5_102 55 149 2.52e-15
R5_11 49 53 0.5
C5_111 49 149 2.4e-15
C5_112 53 149 2.4e-15
R5_12 43 47 0.9
C5_121 43 149 2.52e-15
C5_122 47 149 2.52e-15
R5_13 45 43 0.6
C5_131 45 149 1.75e-15
C5_132 43 149 1.75e-15
R5_14 44 50 650
C5_141 44 149 2.025e-15
C5_142 50 149 2.025e-15
R5_15 46 44 550
C5_151 46 149 1.725e-15
C5_152 44 149 1.725e-15
R4_1 61 64 0.001
R4_2 76 64 0.001
R4_3 62 67 0.001
R4_4 78 67 0.001
R4_5 63 73 0.001
R4_6 79 73 0.001
R4_7 74 75 0.001
C4_71 74 149 2.145e-15
C4_72 75 149 2.145e-15
R4_8 73 74 0.001
C4_81 73 149 2.34e-15
C4_82 74 149 2.34e-15
R4_9 71 73 0.001
C4_91 71 149 1.365e-15
C4_92 73 149 1.365e-15
R4_10 72 71 0.001
C4_101 72 149 3.9e-16
C4_102 71 149 3.9e-16
R4_11 70 72 0.001
C4_111 70 149 1.755e-15
C4_112 72 149 1.755e-15
R4_12 67 70 0.001
C4_121 67 149 2.34e-15
C4_122 70 149 2.34e-15
R4_13 68 67 0.001
C4_131 68 149 1.365e-15
C4_132 67 149 1.365e-15
R4_14 64 66 0.001
C4_141 64 149 2.34e-15
C4_142 66 149 2.34e-15
R4_15 69 68 0.001
C4_151 69 149 3.9e-16
C4_152 68 149 3.9e-16
R4_16 66 69 0.001
C4_161 66 149 1.755e-15
C4_162 69 149 1.755e-15
R4_17 66 77 0.001
C4_171 66 149 7.2e-16
C4_172 77 149 7.2e-16
R4_18 64 77 0.001
C4_181 64 149 7.2e-16
C4_182 77 149 7.2e-16
R4_19 65 64 0.001
C4_191 65 149 1.755e-15
C4_192 64 149 1.755e-15
R3_1 82 83 0.001
R3_2 93 94 0.001
R3_3 102 101 0.001
R3_4 96 95 0.001
R3_5 102 103 0.001
R3_6 98 97 0.001
R3_7 111 110 0.001
R3_8 105 104 0.001
R3_9 90 89 0.001
R3_10 110 112 0.001
R3_11 105 106 0.001
R3_12 108 107 0.001
R3_13 109 118 0.001
R3_14 125 126 0.001
R3_15 114 113 0.001
R3_16 91 92 0.001
R3_17 113 115 0.001
R3_18 117 116 0.001
R3_19 123 124 0.001
R3_20 122 121 0.001
R3_21 122 127 500
C3_211 122 149 1.575e-15
C3_212 127 149 1.575e-15
R3_22 119 122 550
C3_221 119 149 1.65e-15
C3_222 122 149 1.65e-15
R3_23 123 128 500
C3_231 123 149 1.575e-15
C3_232 128 149 1.575e-15
R3_24 120 123 550
C3_241 120 149 1.65e-15
C3_242 123 149 1.65e-15
R3_25 121 130 0.6
C3_251 121 149 1.75e-15
C3_252 130 149 1.75e-15
R3_26 115 121 0.9
C3_261 115 149 2.52e-15
C3_262 121 149 2.52e-15
R3_27 124 131 0.6
C3_271 124 149 1.75e-15
C3_272 131 149 1.75e-15
R3_28 116 124 0.9
C3_281 116 149 2.52e-15
C3_282 124 149 2.52e-15
R3_29 91 100 550
C3_291 91 149 1.65e-15
C3_292 100 149 1.65e-15
R3_30 87 91 500
C3_301 87 149 1.575e-15
C3_302 91 149 1.575e-15
R3_31 113 117 0.35
C3_311 113 149 1.8e-15
C3_312 117 149 1.8e-15
R3_32 92 107 0.9
C3_321 92 149 2.52e-15
C3_322 107 149 2.52e-15
R3_33 88 92 0.6
C3_331 88 149 1.75e-15
C3_332 92 149 1.75e-15
R3_34 106 114 0.5
C3_341 106 149 2.4e-15
C3_342 114 149 2.4e-15
R3_35 126 129 0.001
C3_351 126 149 2.1e-16
C3_352 129 149 2.1e-16
R3_36 118 126 1
C3_361 118 149 2.8e-15
C3_362 126 149 2.8e-15
R3_37 112 118 0.4
C3_371 112 149 1.26e-15
C3_372 118 149 1.26e-15
R3_38 90 99 550
C3_381 90 149 1.65e-15
C3_382 99 149 1.65e-15
R3_39 86 90 500
C3_391 86 149 1.575e-15
C3_392 90 149 1.575e-15
R3_40 105 108 0.35
C3_401 105 149 1.8e-15
C3_402 108 149 1.8e-15
R3_41 97 104 0.2
C3_411 97 149 7e-16
C3_412 104 149 7e-16
R3_42 89 97 0.6
C3_421 89 149 1.82e-15
C3_422 97 149 1.82e-15
R3_43 85 89 0.6
C3_431 85 149 1.75e-15
C3_432 89 149 1.75e-15
R3_44 103 111 0.5
C3_441 103 149 2.4e-15
C3_442 111 149 2.4e-15
R3_45 96 98 0.25
C3_451 96 149 1.2e-15
C3_452 98 149 1.2e-15
R3_46 95 101 0.2
C3_461 95 149 7e-16
C3_462 101 149 7e-16
R3_47 94 95 0.2
C3_471 94 149 5.6e-16
C3_472 95 149 5.6e-16
R3_48 83 94 1
C3_481 83 149 2.8e-15
C3_482 94 149 2.8e-15
R3_49 84 83 0.001
C3_491 84 149 2.1e-16
C3_492 83 149 2.1e-16
R2_1 137 141 0.001
R2_2 142 144 0.001
R2_3 134 135 0.001
R2_4 138 139 0.001
C2_41 138 149 3.6e-16
C2_42 139 149 3.6e-16
R2_5 138 149 0.001
C2_51 138 149 1.2e-15
C2_52 149 149 1.2e-15
R2_6 135 149 0.001
C2_61 135 149 9.6e-16
C2_62 149 149 9.6e-16
R2_7 136 135 0.001
C2_71 136 149 1.08e-15
C2_72 135 149 1.08e-15
R2_8 147 148 0.001
C2_81 147 149 6e-16
C2_82 148 149 6e-16
R2_9 144 147 0.1
C2_91 144 149 2.16e-15
C2_92 147 149 2.16e-15
R2_10 145 144 0.001
C2_101 145 149 8.4e-16
C2_102 144 149 8.4e-16
R2_11 146 145 0.001
C2_111 146 149 2.4e-16
C2_112 145 149 2.4e-16
R2_12 143 146 0.001
C2_121 143 149 3.6e-16
C2_122 146 149 3.6e-16
R2_13 141 143 0.1
C2_131 141 149 2.16e-15
C2_132 143 149 2.16e-15
R2_14 140 141 0.001
C2_141 140 149 8.4e-16
C2_142 141 149 8.4e-16
R2_15 139 140 0.001
C2_151 139 149 2.4e-16
C2_152 140 149 2.4e-16
R1_1 152 153 0.001
R1_2 155 156 0.001
R1_3 156 157 0.4
C1_31 156 149 1.33e-15
C1_32 157 149 1.33e-15
R1_4 153 156 1
C1_41 153 149 2.8e-15
C1_42 156 149 2.8e-15
R1_5 154 153 0.001
C1_51 154 149 2.1e-16
C1_52 153 149 2.1e-16
.ends fo4_gordo2

