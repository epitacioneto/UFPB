* Spice description of noc_roteado
* Spice driver version -1218117063
* Date ( dd/mm/yyyy hh:mm:ss ): 17/11/2020 at 15:44:52

* INTERF ck i10 i5 vdd vss 


.subckt noc_roteado 2 13 10 16 7 
* NET 2 = ck
* NET 3 = i4
* NET 4 = i1
* NET 5 = i2
* NET 6 = i3
* NET 7 = vss
* NET 8 = ck_b
* NET 10 = i5
* NET 11 = i9
* NET 12 = i8
* NET 13 = i10
* NET 14 = i6
* NET 15 = i7
* NET 16 = vdd
Mtr_00026 15 14 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 12 15 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 13 11 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 11 12 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 9 10 14 16 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00021 16 8 9 16 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00020 6 5 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00019 5 4 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00018 3 6 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 1 13 4 16 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00016 16 2 1 16 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00015 10 3 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 8 2 16 16 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00013 7 14 15 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 7 15 12 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 7 11 13 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 7 12 11 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 14 8 7 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 7 10 14 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 7 5 6 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 7 4 5 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 7 6 3 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 4 2 7 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 7 13 4 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00002 7 3 10 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 7 2 8 7 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C15 2 7 5.515e-14
C14 3 7 5.257e-14
C13 4 7 5.481e-14
C12 5 7 5.257e-14
C11 6 7 5.377e-14
C10 7 7 2.3892e-13
C9 8 7 5.114e-14
C7 10 7 5.342e-14
C6 11 7 5.137e-14
C5 12 7 5.497e-14
C4 13 7 5.222e-14
C3 14 7 6.801e-14
C2 15 7 5.017e-14
C1 16 7 2.476e-13
.ends noc_roteado

