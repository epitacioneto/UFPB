
.include inv3_s.spi
* INTERF a vdd vss y1 y2 y3

X1 10 40 30 20 21 22 inv3_s
V1 10 30 dc 0.0V
*RL 20 30 1000k
Vdd 40 30 1.8V
Vss 30 0 0.0V

.model tp pmos level = 54
.model tn nmos level = 54

*.dc V1 0 1.8 0.001
.dc V1 0.716 1.123 0.001
.end
