
.include ff_m_e_noc_roteado.spi
.include latch_d_roteado.spi

* INTERF a ck phi_1 phi_2 q vdd vss 
* INTERF a ck q vdd vss 

X1 20 12 13 14 15 40 30 ff_m_e_noc_roteado
X2 20 12 16 40 30 latch_d_roteado

V1 12 30 pulse(0V 1.8V 50n 1p 1p 50n 100n)
V2 20 30 pulse(0V 1.8V 20n 1p 1p 120n 240n)

*R1 20 0 10Meg 

Vdd 40 0 1.8V
Vss 30 0 0V

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.1ns 960ns
.end
