* Spice description of inversor_equilibrado
* Spice driver version -1218551239
* Date ( dd/mm/yyyy hh:mm:ss ): 17/10/2020 at 20:27:34

* INTERF a vdd vss y 


.subckt inversor_equilibrado 1 13 21 27 
* NET 1 = a
* NET 13 = vdd
* NET 21 = vss
* NET 27 = y
Mtr_00002 30 7 10 13 tp L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00001 26 5 18 21 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R4_1 3 2 0.001
R4_2 1 6 0.7
C4_21 1 21 2.17e-15
C4_22 6 21 2.17e-15
R4_3 2 1 0.1
C4_31 2 21 4.2e-16
C4_32 1 21 4.2e-16
R4_4 4 2 0.6
C4_41 4 21 1.75e-15
C4_42 2 21 1.75e-15
R4_5 3 7 550
C4_51 3 21 1.65e-15
C4_52 7 21 1.65e-15
R4_6 5 3 500
C4_61 5 21 1.575e-15
C4_62 3 21 1.575e-15
R3_1 10 11 0.001
R3_2 14 15 0.001
C3_21 14 21 1.32e-15
C3_22 15 21 1.32e-15
R3_3 14 13 0.001
C3_31 14 21 7.2e-16
C3_32 13 21 7.2e-16
R3_4 11 13 0.001
C3_41 11 21 7.2e-16
C3_42 13 21 7.2e-16
R3_5 12 11 0.001
C3_51 12 21 1.08e-15
C3_52 11 21 1.08e-15
R2_1 18 19 0.001
R2_2 22 23 0.001
C2_21 22 21 6e-16
C2_22 23 21 6e-16
R2_3 22 21 0.001
C2_31 22 21 1.2e-15
C2_32 21 21 1.2e-15
R2_4 19 21 0.001
C2_41 19 21 9.6e-16
C2_42 21 21 9.6e-16
R2_5 20 19 0.001
C2_51 20 21 1.08e-15
C2_52 19 21 1.08e-15
R1_1 26 28 0.001
R1_2 30 31 0.001
R1_3 31 32 0.4
C1_31 31 21 1.33e-15
C1_32 32 21 1.33e-15
R1_4 27 31 0.8
C1_41 27 21 2.24e-15
C1_42 31 21 2.24e-15
R1_5 28 27 0.2
C1_51 28 21 5.6e-16
C1_52 27 21 5.6e-16
R1_6 29 28 0.001
C1_61 29 21 2.1e-16
C1_62 28 21 2.1e-16
.ends inversor_equilibrado

