
.include noc.spi
.include noc_roteado.spi

* INTERF phi phi1 phi2 vdd vss vss1 
* INTERF ck i10 i5 vdd vss

X1 20 10 11 40 30 30 noc
X2 20 12 13 40 30 noc_roteado

V1 20 0 pulse(0V 1.8V 7n 1p 1p 5n 10n)

*R1 20 0 10Meg 

Vdd 40 0 1.8V
Vss 30 0 0V

.model tp pmos level = 54
.model tn nmos level = 54

.tran 0.01ns 40ns
.end
