* Spice description of trans_gate
* Spice driver version -1218551239
* Date ( dd/mm/yyyy hh:mm:ss ):  3/11/2020 at 15:05:46

* INTERF a enable vdd vss y 


.subckt trans_gate 58 9 14 35 50 
* NET 9 = enable
* NET 14 = vdd
* NET 35 = vss
* NET 50 = y
* NET 58 = a
Mtr_00004 59 28 49 14 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 26 6 13 14 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 55 4 45 35 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 23 1 36 35 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R6_1 8 7 0.001
R6_2 9 10 0.2
C6_21 9 35 7.7e-16
C6_22 10 35 7.7e-16
R6_3 7 9 0.6
C6_31 7 35 1.82e-15
C6_32 9 35 1.82e-15
R6_4 2 7 0.6
C6_41 2 35 1.75e-15
C6_42 7 35 1.75e-15
R6_5 8 6 450
C6_51 8 35 1.425e-15
C6_52 6 35 1.425e-15
R6_6 1 8 500
C6_61 1 35 1.575e-15
C6_62 8 35 1.575e-15
R6_7 3 1 150
C6_71 3 35 5.25e-16
C6_72 1 35 5.25e-16
R6_8 3 5 800
C6_81 3 35 2.4e-15
C6_82 5 35 2.4e-15
R6_9 5 4 150
C6_91 5 35 5.25e-16
C6_92 4 35 5.25e-16
R5_1 13 14 0.001
R5_2 19 18 0.001
R5_3 18 20 0.001
C5_31 18 35 1.08e-15
C5_32 20 35 1.08e-15
R5_4 16 18 0.1
C5_41 16 35 2.52e-15
C5_42 18 35 2.52e-15
R5_5 17 16 0.001
C5_51 17 35 2.4e-16
C5_52 16 35 2.4e-16
R5_6 14 17 0.1
C5_61 14 35 2.52e-15
C5_62 17 35 2.52e-15
R5_7 15 14 0.001
C5_71 15 35 1.08e-15
C5_72 14 35 1.08e-15
R4_1 23 24 0.001
R4_2 30 29 0.001
R4_3 26 27 0.001
R4_4 28 31 300
C4_41 28 35 9.75e-16
C4_42 31 35 9.75e-16
R4_5 30 31 650
C4_51 30 35 1.95e-15
C4_52 31 35 1.95e-15
R4_6 29 32 0.1
C4_61 29 35 3.5e-16
C4_62 32 35 3.5e-16
R4_7 27 29 0.3
C4_71 27 35 9.8e-16
C4_72 29 35 9.8e-16
R4_8 24 27 1
C4_81 24 35 2.8e-15
C4_82 27 35 2.8e-15
R4_9 25 24 0.001
C4_91 25 35 2.1e-16
C4_92 24 35 2.1e-16
R3_1 36 35 0.001
R3_2 41 40 0.001
R3_3 40 42 0.001
C3_31 40 35 1.08e-15
C3_32 42 35 1.08e-15
R3_4 38 40 0.1
C3_41 38 35 2.52e-15
C3_42 40 35 2.52e-15
R3_5 39 38 0.001
C3_51 39 35 2.4e-16
C3_52 38 35 2.4e-16
R3_6 35 39 0.1
C3_61 35 35 2.52e-15
C3_62 39 35 2.52e-15
R3_7 37 35 0.001
C3_71 37 35 1.08e-15
C3_72 35 35 1.08e-15
R2_1 45 46 0.001
R2_2 49 51 0.001
R2_3 51 52 0.1
C2_31 51 35 1.725e-16
C2_32 52 35 1.725e-16
R2_4 50 51 0.3
C2_41 50 35 3.45e-16
C2_42 51 35 3.45e-16
R2_5 47 50 1.3
C2_51 47 35 1.5525e-15
C2_52 50 35 1.5525e-15
R2_6 48 47 0.2
C2_61 48 35 2.3e-16
C2_62 47 35 2.3e-16
R2_7 46 48 0.1
C2_71 46 35 1.725e-16
C2_72 48 35 1.725e-16
R1_1 55 56 0.001
R1_2 59 60 0.001
R1_3 60 61 0.4
C1_31 60 35 1.33e-15
C1_32 61 35 1.33e-15
R1_4 58 60 0.3
C1_41 58 35 8.4e-16
C1_42 60 35 8.4e-16
R1_5 56 58 0.7
C1_51 56 35 1.96e-15
C1_52 58 35 1.96e-15
R1_6 57 56 0.001
C1_61 57 35 2.1e-16
C1_62 56 35 2.1e-16
.ends trans_gate

