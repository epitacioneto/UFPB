* Spice description of mux_4_n_inverter
* Spice driver version -1217678791
* Date ( dd/mm/yyyy hh:mm:ss ): 10/11/2020 at 16:10:26

* INTERF d0 d1 d2 d3 s0 s1 vdd vss vss1 y 


.subckt mux_4_n_inverter 43 34 110 52 86 223 300 356 31 346 
* NET 31 = vss1
* NET 34 = d1
* NET 43 = d0
* NET 52 = d3
* NET 86 = s0
* NET 110 = d2
* NET 223 = s1
* NET 300 = vdd
* NET 346 = y
* NET 356 = vss
Mtr_00028 293 206 347 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00027 293 260 296 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00026 290 241 349 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00025 290 190 297 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00024 163 75 191 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00023 163 116 298 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00022 61 126 193 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00021 61 58 299 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00020 7 91 266 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00019 7 45 327 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00018 1 147 269 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00017 1 36 328 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00016 139 87 326 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00015 250 219 325 300 tp L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00014 373 230 336 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00013 373 257 355 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00012 333 205 341 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00011 333 169 358 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00010 166 122 171 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00009 166 114 362 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00008 64 67 174 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00007 64 56 366 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00006 10 159 274 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00005 10 49 15 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00004 4 106 283 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00003 4 40 16 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00002 152 104 14 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
Mtr_00001 252 226 13 356 tn L=1U W=2U AS=4P AD=4P PS=8U PD=8U 
R22_1 13 17 0.001
R22_2 14 21 0.001
R22_3 15 24 0.001
R22_4 16 27 0.001
R22_5 27 30 0.2
C22_51 27 356 3.96e-15
C22_52 30 356 3.96e-15
R22_6 28 27 0.001
C22_61 28 356 8.4e-16
C22_62 27 356 8.4e-16
R22_7 29 28 0.001
C22_71 29 356 2.4e-16
C22_72 28 356 2.4e-16
R22_8 24 29 0.2
C22_81 24 356 3.72e-15
C22_82 29 356 3.72e-15
R22_9 25 24 0.001
C22_91 25 356 8.4e-16
C22_92 24 356 8.4e-16
R22_10 26 25 0.001
C22_101 26 356 2.4e-16
C22_102 25 356 2.4e-16
R22_11 20 26 0.001
C22_111 20 356 3.6e-16
C22_112 26 356 3.6e-16
R22_12 21 20 0.1
C22_121 21 356 2.16e-15
C22_122 20 356 2.16e-15
R22_13 22 21 0.001
C22_131 22 356 8.4e-16
C22_132 21 356 8.4e-16
R22_14 23 22 0.001
C22_141 23 356 2.4e-16
C22_142 22 356 2.4e-16
R22_15 17 23 0.001
C22_151 17 356 8.4e-16
C22_152 23 356 8.4e-16
R22_16 17 31 0.001
C22_161 17 356 9.6e-16
C22_162 31 356 9.6e-16
R22_17 18 31 0.001
C22_171 18 356 1.2e-15
C22_172 31 356 1.2e-15
R22_18 19 18 0.001
C22_181 19 356 6e-16
C22_182 18 356 6e-16
R21_1 38 37 0.001
R21_2 38 40 500
C21_21 38 356 1.575e-15
C21_22 40 356 1.575e-15
R21_3 36 38 450
C21_31 36 356 1.425e-15
C21_32 38 356 1.425e-15
R21_4 37 39 0.6
C21_41 37 356 1.75e-15
C21_42 39 356 1.75e-15
R21_5 34 37 0.1
C21_51 34 356 4.2e-16
C21_52 37 356 4.2e-16
R21_6 35 34 0.7
C21_61 35 356 2.17e-15
C21_62 34 356 2.17e-15
R20_1 47 46 0.001
R20_2 47 49 500
C20_21 47 356 1.575e-15
C20_22 49 356 1.575e-15
R20_3 45 47 450
C20_31 45 356 1.425e-15
C20_32 47 356 1.425e-15
R20_4 46 48 0.6
C20_41 46 356 1.75e-15
C20_42 48 356 1.75e-15
R20_5 43 46 0.1
C20_51 43 356 4.2e-16
C20_52 46 356 4.2e-16
R20_6 44 43 0.7
C20_61 44 356 2.17e-15
C20_62 43 356 2.17e-15
R19_1 54 53 0.001
R19_2 52 57 0.7
C19_21 52 356 2.17e-15
C19_22 57 356 2.17e-15
R19_3 53 52 0.1
C19_31 53 356 4.2e-16
C19_32 52 356 4.2e-16
R19_4 55 53 0.6
C19_41 55 356 1.75e-15
C19_42 53 356 1.75e-15
R19_5 54 58 450
C19_51 54 356 1.425e-15
C19_52 58 356 1.425e-15
R19_6 56 54 500
C19_61 56 356 1.575e-15
C19_62 54 356 1.575e-15
R16_1 80 79 0.001
R16_2 74 73 0.001
R16_3 77 76 0.001
R16_4 93 92 0.001
R16_5 69 68 0.001
R16_6 99 98 0.001
R16_7 101 100 0.001
R16_8 68 70 0.001
R16_9 89 88 0.001
R16_10 100 102 0.001
R16_11 95 94 0.001
R16_12 70 71 0.001
R16_13 102 103 0.001
R16_14 85 84 0.001
R16_15 97 96 0.001
R16_16 103 106 400
C16_161 103 356 1.275e-15
C16_162 106 356 1.275e-15
R16_17 96 104 500
C16_171 96 356 1.575e-15
C16_172 104 356 1.575e-15
R16_18 87 96 450
C16_181 87 356 1.425e-15
C16_182 96 356 1.425e-15
R16_19 85 91 350
C16_191 85 356 1.125e-15
C16_192 91 356 1.125e-15
R16_20 67 71 400
C16_201 67 356 1.275e-15
C16_202 71 356 1.275e-15
R16_21 102 107 1
C16_211 102 356 1.2075e-15
C16_212 107 356 1.2075e-15
R16_22 97 105 0.6
C16_221 97 356 1.75e-15
C16_222 105 356 1.75e-15
R16_23 94 97 0.1
C16_231 94 356 4.2e-16
C16_232 97 356 4.2e-16
R16_24 86 94 0.2
C16_241 86 356 7e-16
C16_242 94 356 7e-16
R16_25 82 86 0.5
C16_251 82 356 1.47e-15
C16_252 86 356 1.47e-15
R16_26 90 84 0.5
C16_261 90 356 5.75e-16
C16_262 84 356 5.75e-16
R16_27 72 70 1
C16_271 72 356 1.2075e-15
C16_272 70 356 1.2075e-15
R16_28 90 88 0.9
C16_281 90 356 1.035e-15
C16_282 88 356 1.035e-15
R16_29 83 90 0.2
C16_291 83 356 2.875e-16
C16_292 90 356 2.875e-16
R16_30 95 98 1
C16_301 95 356 4.8e-15
C16_302 98 356 4.8e-15
R16_31 89 92 0.5
C16_311 89 356 2.4e-15
C16_312 92 356 2.4e-15
R16_32 99 101 0.1
C16_321 99 356 6e-16
C16_322 101 356 6e-16
R16_33 93 99 0.1
C16_331 93 356 6e-16
C16_332 99 356 6e-16
R16_34 69 77 0.25
C16_341 69 356 1.2e-15
C16_342 77 356 1.2e-15
R16_35 77 93 1
C16_351 77 356 4.8e-15
C16_352 93 356 4.8e-15
R16_36 74 76 0.5
C16_361 74 356 2.4e-15
C16_362 76 356 2.4e-15
R16_37 78 81 0.2
C16_371 78 356 2.875e-16
C16_372 81 356 2.875e-16
R16_38 73 78 0.9
C16_381 73 356 1.035e-15
C16_382 78 356 1.035e-15
R16_39 78 79 0.5
C16_391 78 356 5.75e-16
C16_392 79 356 5.75e-16
R16_40 75 80 350
C16_401 75 356 1.125e-15
C16_402 80 356 1.125e-15
R15_1 112 111 0.001
R15_2 110 115 0.7
C15_21 110 356 2.17e-15
C15_22 115 356 2.17e-15
R15_3 111 110 0.1
C15_31 111 356 4.2e-16
C15_32 110 356 4.2e-16
R15_4 113 111 0.6
C15_41 113 356 1.75e-15
C15_42 111 356 1.75e-15
R15_5 112 116 450
C15_51 112 356 1.425e-15
C15_52 116 356 1.425e-15
R15_6 114 112 500
C15_61 114 356 1.575e-15
C15_62 112 356 1.575e-15
R14_1 123 119 0.001
R14_2 119 120 0.001
R14_3 120 121 0.001
R14_4 128 127 0.001
R14_5 142 141 0.001
R14_6 130 129 0.001
R14_7 149 148 0.001
R14_8 144 143 0.001
R14_9 148 150 0.001
R14_10 133 132 0.001
R14_11 150 151 0.001
R14_12 138 137 0.001
R14_13 158 157 0.001
R14_14 154 153 0.001
R14_15 139 140 0.001
R14_16 152 155 0.001
R14_17 155 156 0.001
C14_171 155 356 2.1e-16
C14_172 156 356 2.1e-16
R14_18 153 155 0.2
C14_181 153 356 5.6e-16
C14_182 155 356 5.6e-16
R14_19 140 153 0.8
C14_191 140 356 2.24e-15
C14_192 153 356 2.24e-15
R14_20 135 140 0.4
C14_201 135 356 1.33e-15
C14_202 140 356 1.33e-15
R14_21 151 159 400
C14_211 151 356 1.275e-15
C14_212 159 356 1.275e-15
R14_22 138 147 350
C14_221 138 356 1.125e-15
C14_222 147 356 1.125e-15
R14_23 154 158 0.35
C14_231 154 356 1.8e-15
C14_232 158 356 1.8e-15
R14_24 126 133 350
C14_241 126 356 1.125e-15
C14_242 133 356 1.125e-15
R14_25 157 160 0.5
C14_251 157 356 6.325e-16
C14_252 160 356 6.325e-16
R14_26 150 157 0.5
C14_261 150 356 5.75e-16
C14_262 157 356 5.75e-16
R14_27 145 137 0.5
C14_271 145 356 5.75e-16
C14_272 137 356 5.75e-16
R14_28 143 146 0.5
C14_281 143 356 6.325e-16
C14_282 146 356 6.325e-16
R14_29 145 143 0.4
C14_291 145 356 4.6e-16
C14_292 143 356 4.6e-16
R14_30 136 145 0.2
C14_301 136 356 2.875e-16
C14_302 145 356 2.875e-16
R14_31 131 132 0.5
C14_311 131 356 5.75e-16
C14_312 132 356 5.75e-16
R14_32 131 134 0.2
C14_321 131 356 2.875e-16
C14_322 134 356 2.875e-16
R14_33 129 131 0.4
C14_331 129 356 4.6e-16
C14_332 131 356 4.6e-16
R14_34 125 129 0.5
C14_341 125 356 6.325e-16
C14_342 129 356 6.325e-16
R14_35 141 144 0.5
C14_351 141 356 2.4e-15
C14_352 144 356 2.4e-15
R14_36 142 149 0.35
C14_361 142 356 1.8e-15
C14_362 149 356 1.8e-15
R14_37 127 130 0.5
C14_371 127 356 2.4e-15
C14_372 130 356 2.4e-15
R14_38 128 142 0.75
C14_381 128 356 3.6e-15
C14_382 142 356 3.6e-15
R14_39 121 128 0.35
C14_391 121 356 1.8e-15
C14_392 128 356 1.8e-15
R14_40 124 119 1
C14_401 124 356 1.2075e-15
C14_402 119 356 1.2075e-15
R14_41 122 123 400
C14_411 122 356 1.275e-15
C14_412 123 356 1.275e-15
R11_1 182 181 0.001
R11_2 183 181 0.001
R11_3 183 184 0.001
R11_4 184 185 0.001
R11_5 187 186 0.001
R11_6 186 188 0.001
R11_7 188 189 0.001
R11_8 191 192 0.001
R11_9 178 177 0.001
R11_10 171 172 0.001
R11_11 180 179 0.001
R11_12 193 194 0.001
R11_13 174 175 0.001
R11_14 175 176 0.1
C11_141 175 356 1.725e-16
C11_142 176 356 1.725e-16
R11_15 194 196 0.1
C11_151 194 356 1.725e-16
C11_152 196 356 1.725e-16
R11_16 179 194 1.6
C11_161 179 356 1.84e-15
C11_162 194 356 1.84e-15
R11_17 176 179 0.2
C11_171 176 356 2.875e-16
C11_172 179 356 2.875e-16
R11_18 178 180 0.5
C11_181 178 356 2.4e-15
C11_182 180 356 2.4e-15
R11_19 172 173 0.1
C11_191 172 356 1.725e-16
C11_192 173 356 1.725e-16
R11_20 192 195 0.1
C11_201 192 356 1.725e-16
C11_202 195 356 1.725e-16
R11_21 189 192 1.1
C11_211 189 356 1.265e-15
C11_212 192 356 1.265e-15
R11_22 177 189 0.5
C11_221 177 356 5.75e-16
C11_222 189 356 5.75e-16
R11_23 173 177 0.2
C11_231 173 356 2.875e-16
C11_232 177 356 2.875e-16
R11_24 185 187 0.75
C11_241 185 356 3.72e-15
C11_242 187 356 3.72e-15
R11_25 181 197 0.9
C11_251 181 356 2.73e-15
C11_252 197 356 2.73e-15
R11_26 170 181 0.5
C11_261 170 356 1.61e-15
C11_262 181 356 1.61e-15
R11_27 182 190 450
C11_271 182 356 1.425e-15
C11_272 190 356 1.425e-15
R11_28 169 182 500
C11_281 169 356 1.575e-15
C11_282 182 356 1.575e-15
R10_1 215 218 0.001
R10_2 208 207 0.001
R10_3 212 211 0.001
R10_4 214 213 0.001
R10_5 201 200 0.001
R10_6 200 202 0.001
R10_7 210 209 0.001
R10_8 202 203 0.001
R10_9 221 220 0.001
R10_10 220 222 0.001
R10_11 225 224 0.001
R10_12 225 226 500
C10_121 225 356 1.575e-15
C10_122 226 356 1.575e-15
R10_13 219 225 450
C10_131 219 356 1.425e-15
C10_132 225 356 1.425e-15
R10_14 224 227 0.6
C10_141 224 356 1.75e-15
C10_142 227 356 1.75e-15
R10_15 223 224 0.1
C10_151 223 356 4.2e-16
C10_152 224 356 4.2e-16
R10_16 222 223 0.7
C10_161 222 356 2.1e-15
C10_162 223 356 2.1e-15
R10_17 205 203 400
C10_171 205 356 1.275e-15
C10_172 203 356 1.275e-15
R10_18 204 202 1
C10_181 204 356 1.2075e-15
C10_182 202 356 1.2075e-15
R10_19 210 221 0.85
C10_191 210 356 4.2e-15
C10_192 221 356 4.2e-15
R10_20 209 213 0.25
C10_201 209 356 1.2e-15
C10_202 213 356 1.2e-15
R10_21 214 211 0.1
C10_211 214 356 6e-16
C10_212 211 356 6e-16
R10_22 201 214 0.1
C10_221 201 356 6e-16
C10_222 214 356 6e-16
R10_23 208 212 0.5
C10_231 208 356 2.4e-15
C10_232 212 356 2.4e-15
R10_24 216 217 0.2
C10_241 216 356 2.875e-16
C10_242 217 356 2.875e-16
R10_25 207 216 0.9
C10_251 207 356 1.035e-15
C10_252 216 356 1.035e-15
R10_26 216 218 0.5
C10_261 216 356 5.75e-16
C10_262 218 356 5.75e-16
R10_27 206 215 350
C10_271 206 356 1.125e-15
C10_272 215 356 1.125e-15
R9_1 232 231 0.001
R9_2 231 233 0.001
R9_3 233 234 0.001
R9_4 237 236 0.001
R9_5 247 246 0.001
R9_6 239 238 0.001
R9_7 249 248 0.001
R9_8 245 244 0.001
R9_9 250 251 0.001
R9_10 252 253 0.001
R9_11 241 245 350
C9_111 241 356 1.125e-15
C9_112 245 356 1.125e-15
R9_12 253 254 0.001
C9_121 253 356 2.1e-16
C9_122 254 356 2.1e-16
R9_13 251 253 1
C9_131 251 356 2.8e-15
C9_132 253 356 2.8e-15
R9_14 248 251 0.4
C9_141 248 356 1.26e-15
C9_142 251 356 1.26e-15
R9_15 242 244 0.5
C9_151 242 356 5.75e-16
C9_152 244 356 5.75e-16
R9_16 242 243 0.2
C9_161 242 356 2.875e-16
C9_162 243 356 2.875e-16
R9_17 238 242 0.4
C9_171 238 356 4.6e-16
C9_172 242 356 4.6e-16
R9_18 240 238 0.5
C9_181 240 356 6.325e-16
C9_182 238 356 6.325e-16
R9_19 246 249 0.1
C9_191 246 356 6e-16
C9_192 249 356 6e-16
R9_20 236 239 0.5
C9_201 236 356 2.4e-15
C9_202 239 356 2.4e-15
R9_21 237 247 0.6
C9_211 237 356 3e-15
C9_212 247 356 3e-15
R9_22 234 237 0.35
C9_221 234 356 1.8e-15
C9_222 237 356 1.8e-15
R9_23 235 231 1
C9_231 235 356 1.2075e-15
C9_232 231 356 1.2075e-15
R9_24 230 232 400
C9_241 230 356 1.275e-15
C9_242 232 356 1.275e-15
R8_1 258 261 0.001
R8_2 263 262 0.001
R8_3 263 264 0.001
R8_4 264 265 0.001
R8_5 273 272 0.001
R8_6 276 275 0.001
R8_7 275 277 0.001
R8_8 277 278 0.001
R8_9 266 267 0.001
R8_10 280 279 0.001
R8_11 274 281 0.001
R8_12 285 284 0.001
R8_13 269 270 0.001
R8_14 283 286 0.001
R8_15 287 286 0.1
C8_151 287 356 1.725e-16
C8_152 286 356 1.725e-16
R8_16 284 287 0.2
C8_161 284 356 2.875e-16
C8_162 287 356 2.875e-16
R8_17 270 284 1.6
C8_171 270 356 1.84e-15
C8_172 284 356 1.84e-15
R8_18 271 270 0.1
C8_181 271 356 1.725e-16
C8_182 270 356 1.725e-16
R8_19 280 285 0.5
C8_191 280 356 2.4e-15
C8_192 285 356 2.4e-15
R8_20 282 281 0.1
C8_201 282 356 1.725e-16
C8_202 281 356 1.725e-16
R8_21 279 282 0.2
C8_211 279 356 2.875e-16
C8_212 282 356 2.875e-16
R8_22 278 279 0.5
C8_221 278 356 5.75e-16
C8_222 279 356 5.75e-16
R8_23 267 278 1.1
C8_231 267 356 1.265e-15
C8_232 278 356 1.265e-15
R8_24 268 267 0.1
C8_241 268 356 1.725e-16
C8_242 267 356 1.725e-16
R8_25 273 276 1.3
C8_251 273 356 6.24e-15
C8_252 276 356 6.24e-15
R8_26 264 272 1
C8_261 264 356 4.8e-15
C8_262 272 356 4.8e-15
R8_27 261 262 0.9
C8_271 261 356 2.52e-15
C8_272 262 356 2.52e-15
R8_28 259 261 0.6
C8_281 259 356 1.75e-15
C8_282 261 356 1.75e-15
R8_29 258 260 450
C8_291 258 356 1.425e-15
C8_292 260 356 1.425e-15
R8_30 257 258 500
C8_301 257 356 1.575e-15
C8_302 258 356 1.575e-15
R5_1 296 300 0.001
R5_2 304 303 0.001
R5_3 310 309 0.001
R5_4 297 305 0.001
R5_5 325 306 0.001
R5_6 298 312 0.001
R5_7 317 316 0.001
R5_8 327 312 0.001
R5_9 329 316 0.001
R5_10 326 311 0.001
R5_11 328 321 0.001
R5_12 330 322 0.001
R5_13 299 321 0.001
R5_14 323 322 0.001
R5_15 322 324 0.001
C5_151 322 356 1.755e-15
C5_152 324 356 1.755e-15
R5_16 320 322 0.001
C5_161 320 356 2.34e-15
C5_162 322 356 2.34e-15
R5_17 321 320 0.001
C5_171 321 356 2.34e-15
C5_172 320 356 2.34e-15
R5_18 318 321 0.001
C5_181 318 356 1.365e-15
C5_182 321 356 1.365e-15
R5_19 319 318 0.001
C5_191 319 356 3.9e-16
C5_192 318 356 3.9e-16
R5_20 316 319 0.001
C5_201 316 356 1.365e-15
C5_202 319 356 1.365e-15
R5_21 315 316 0.001
C5_211 315 356 2.34e-15
C5_212 316 356 2.34e-15
R5_22 312 315 0.001
C5_221 312 356 2.34e-15
C5_222 315 356 2.34e-15
R5_23 314 312 0.001
C5_231 314 356 1.365e-15
C5_232 312 356 1.365e-15
R5_24 313 314 0.001
C5_241 313 356 3.9e-16
C5_242 314 356 3.9e-16
R5_25 309 313 0.001
C5_251 309 356 1.56e-15
C5_252 313 356 1.56e-15
R5_26 311 309 0.001
C5_261 311 356 2.34e-15
C5_262 309 356 2.34e-15
R5_27 307 311 0.001
C5_271 307 356 1.56e-15
C5_272 311 356 1.56e-15
R5_28 305 307 0.001
C5_281 305 356 5.85e-16
C5_282 307 356 5.85e-16
R5_29 306 305 0.001
C5_291 306 356 1.17e-15
C5_292 305 356 1.17e-15
R5_30 308 306 0.001
C5_301 308 356 5.85e-16
C5_302 306 356 5.85e-16
R5_31 303 308 0.001
C5_311 303 356 1.56e-15
C5_312 308 356 1.56e-15
R5_32 302 303 0.001
C5_321 302 356 2.145e-15
C5_322 303 356 2.145e-15
R5_33 300 302 0.1
C5_331 300 356 1.44e-15
C5_332 302 356 1.44e-15
R5_34 301 300 0.001
C5_341 301 356 1.08e-15
C5_342 300 356 1.08e-15
R3_1 336 337 0.001
R3_2 339 338 0.001
R3_3 347 348 0.001
R3_4 343 342 0.001
R3_5 341 344 0.001
R3_6 349 350 0.001
R3_7 350 352 0.1
C3_71 350 356 1.725e-16
C3_72 352 356 1.725e-16
R3_8 346 350 0.6
C3_81 346 356 6.9e-16
C3_82 350 356 6.9e-16
R3_9 342 346 1
C3_91 342 356 1.15e-15
C3_92 346 356 1.15e-15
R3_10 345 342 0.2
C3_101 345 356 2.875e-16
C3_102 342 356 2.875e-16
R3_11 344 345 0.1
C3_111 344 356 1.725e-16
C3_112 345 356 1.725e-16
R3_12 339 343 0.5
C3_121 339 356 2.4e-15
C3_122 343 356 2.4e-15
R3_13 348 351 0.1
C3_131 348 356 1.725e-16
C3_132 351 356 1.725e-16
R3_14 338 348 1.6
C3_141 338 356 1.84e-15
C3_142 348 356 1.84e-15
R3_15 340 338 0.2
C3_151 340 356 2.875e-16
C3_152 338 356 2.875e-16
R3_16 337 340 0.1
C3_161 337 356 1.725e-16
C3_162 340 356 1.725e-16
R2_1 355 356 0.001
R2_2 358 359 0.001
R2_3 362 363 0.001
R2_4 366 367 0.001
R2_5 367 370 0.2
C2_51 367 356 3.96e-15
C2_52 370 356 3.96e-15
R2_6 368 367 0.001
C2_61 368 356 8.4e-16
C2_62 367 356 8.4e-16
R2_7 369 368 0.001
C2_71 369 356 2.4e-16
C2_72 368 356 2.4e-16
R2_8 363 369 0.2
C2_81 363 356 3.72e-15
C2_82 369 356 3.72e-15
R2_9 364 363 0.001
C2_91 364 356 8.4e-16
C2_92 363 356 8.4e-16
R2_10 365 364 0.001
C2_101 365 356 2.4e-16
C2_102 364 356 2.4e-16
R2_11 359 365 0.2
C2_111 359 356 3.72e-15
C2_112 365 356 3.72e-15
R2_12 360 359 0.001
C2_121 360 356 8.4e-16
C2_122 359 356 8.4e-16
R2_13 361 360 0.001
C2_131 361 356 2.4e-16
C2_132 360 356 2.4e-16
R2_14 356 361 0.2
C2_141 356 356 3.72e-15
C2_142 361 356 3.72e-15
R2_15 357 356 0.001
C2_151 357 356 1.08e-15
C2_152 356 356 1.08e-15
.ends mux_4_n_inverter

