
.include tran_passagem.spi

* INTERF a enable vdd vss y1 y2 

X1 10 11 40 30 20 21 tran_passagem
V1 10 0 dc 0.0V
V2 11 0 dc 1.8V

R1 21 0 100k
R2 20 0 100k 

Vdd 40 0 1.8V
Vss 30 0 -1.8V

.model tp pmos level = 54
.model tn nmos level = 54

.dc V1 -1.8 1.8 0.001
.end

